
// 	Tue Jan  3 00:12:11 2023
//	vlsi
//	localhost.localdomain

module datapath__0_12 (multiplicand, accumulator, p_0);

output [63:0] p_0;
input [63:0] accumulator;
input [63:0] multiplicand;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;


XNOR2_X1 i_64 (.ZN (p_0[63]), .A (n_63), .B (n_62));
XNOR2_X1 i_63 (.ZN (n_63), .A (multiplicand[63]), .B (accumulator[63]));
FA_X1 i_62 (.CO (n_62), .S (p_0[62]), .A (multiplicand[62]), .B (accumulator[62]), .CI (n_61));
FA_X1 i_61 (.CO (n_61), .S (p_0[61]), .A (multiplicand[61]), .B (accumulator[61]), .CI (n_60));
FA_X1 i_60 (.CO (n_60), .S (p_0[60]), .A (multiplicand[60]), .B (accumulator[60]), .CI (n_59));
FA_X1 i_59 (.CO (n_59), .S (p_0[59]), .A (multiplicand[59]), .B (accumulator[59]), .CI (n_58));
FA_X1 i_58 (.CO (n_58), .S (p_0[58]), .A (multiplicand[58]), .B (accumulator[58]), .CI (n_57));
FA_X1 i_57 (.CO (n_57), .S (p_0[57]), .A (multiplicand[57]), .B (accumulator[57]), .CI (n_56));
FA_X1 i_56 (.CO (n_56), .S (p_0[56]), .A (multiplicand[56]), .B (accumulator[56]), .CI (n_55));
FA_X1 i_55 (.CO (n_55), .S (p_0[55]), .A (multiplicand[55]), .B (accumulator[55]), .CI (n_54));
FA_X1 i_54 (.CO (n_54), .S (p_0[54]), .A (multiplicand[54]), .B (accumulator[54]), .CI (n_53));
FA_X1 i_53 (.CO (n_53), .S (p_0[53]), .A (multiplicand[53]), .B (accumulator[53]), .CI (n_52));
FA_X1 i_52 (.CO (n_52), .S (p_0[52]), .A (multiplicand[52]), .B (accumulator[52]), .CI (n_51));
FA_X1 i_51 (.CO (n_51), .S (p_0[51]), .A (multiplicand[51]), .B (accumulator[51]), .CI (n_50));
FA_X1 i_50 (.CO (n_50), .S (p_0[50]), .A (multiplicand[50]), .B (accumulator[50]), .CI (n_49));
FA_X1 i_49 (.CO (n_49), .S (p_0[49]), .A (multiplicand[49]), .B (accumulator[49]), .CI (n_48));
FA_X1 i_48 (.CO (n_48), .S (p_0[48]), .A (multiplicand[48]), .B (accumulator[48]), .CI (n_47));
FA_X1 i_47 (.CO (n_47), .S (p_0[47]), .A (multiplicand[47]), .B (accumulator[47]), .CI (n_46));
FA_X1 i_46 (.CO (n_46), .S (p_0[46]), .A (multiplicand[46]), .B (accumulator[46]), .CI (n_45));
FA_X1 i_45 (.CO (n_45), .S (p_0[45]), .A (multiplicand[45]), .B (accumulator[45]), .CI (n_44));
FA_X1 i_44 (.CO (n_44), .S (p_0[44]), .A (multiplicand[44]), .B (accumulator[44]), .CI (n_43));
FA_X1 i_43 (.CO (n_43), .S (p_0[43]), .A (multiplicand[43]), .B (accumulator[43]), .CI (n_42));
FA_X1 i_42 (.CO (n_42), .S (p_0[42]), .A (multiplicand[42]), .B (accumulator[42]), .CI (n_41));
FA_X1 i_41 (.CO (n_41), .S (p_0[41]), .A (multiplicand[41]), .B (accumulator[41]), .CI (n_40));
FA_X1 i_40 (.CO (n_40), .S (p_0[40]), .A (multiplicand[40]), .B (accumulator[40]), .CI (n_39));
FA_X1 i_39 (.CO (n_39), .S (p_0[39]), .A (multiplicand[39]), .B (accumulator[39]), .CI (n_38));
FA_X1 i_38 (.CO (n_38), .S (p_0[38]), .A (multiplicand[38]), .B (accumulator[38]), .CI (n_37));
FA_X1 i_37 (.CO (n_37), .S (p_0[37]), .A (multiplicand[37]), .B (accumulator[37]), .CI (n_36));
FA_X1 i_36 (.CO (n_36), .S (p_0[36]), .A (multiplicand[36]), .B (accumulator[36]), .CI (n_35));
FA_X1 i_35 (.CO (n_35), .S (p_0[35]), .A (multiplicand[35]), .B (accumulator[35]), .CI (n_34));
FA_X1 i_34 (.CO (n_34), .S (p_0[34]), .A (multiplicand[34]), .B (accumulator[34]), .CI (n_33));
FA_X1 i_33 (.CO (n_33), .S (p_0[33]), .A (multiplicand[33]), .B (accumulator[33]), .CI (n_32));
FA_X1 i_32 (.CO (n_32), .S (p_0[32]), .A (multiplicand[32]), .B (accumulator[32]), .CI (n_31));
FA_X1 i_31 (.CO (n_31), .S (p_0[31]), .A (multiplicand[31]), .B (accumulator[31]), .CI (n_30));
FA_X1 i_30 (.CO (n_30), .S (p_0[30]), .A (multiplicand[30]), .B (accumulator[30]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (p_0[29]), .A (multiplicand[29]), .B (accumulator[29]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (p_0[28]), .A (multiplicand[28]), .B (accumulator[28]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (p_0[27]), .A (multiplicand[27]), .B (accumulator[27]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (p_0[26]), .A (multiplicand[26]), .B (accumulator[26]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (p_0[25]), .A (multiplicand[25]), .B (accumulator[25]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (p_0[24]), .A (multiplicand[24]), .B (accumulator[24]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (p_0[23]), .A (multiplicand[23]), .B (accumulator[23]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (p_0[22]), .A (multiplicand[22]), .B (accumulator[22]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (p_0[21]), .A (multiplicand[21]), .B (accumulator[21]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (p_0[20]), .A (multiplicand[20]), .B (accumulator[20]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (p_0[19]), .A (multiplicand[19]), .B (accumulator[19]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (p_0[18]), .A (multiplicand[18]), .B (accumulator[18]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (p_0[17]), .A (multiplicand[17]), .B (accumulator[17]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (p_0[16]), .A (multiplicand[16]), .B (accumulator[16]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (p_0[15]), .A (multiplicand[15]), .B (accumulator[15]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (p_0[14]), .A (multiplicand[14]), .B (accumulator[14]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (p_0[13]), .A (multiplicand[13]), .B (accumulator[13]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (p_0[12]), .A (multiplicand[12]), .B (accumulator[12]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (p_0[11]), .A (multiplicand[11]), .B (accumulator[11]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (p_0[10]), .A (multiplicand[10]), .B (accumulator[10]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (p_0[9]), .A (multiplicand[9]), .B (accumulator[9]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (p_0[8]), .A (multiplicand[8]), .B (accumulator[8]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (p_0[7]), .A (multiplicand[7]), .B (accumulator[7]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (p_0[6]), .A (multiplicand[6]), .B (accumulator[6]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (p_0[5]), .A (multiplicand[5]), .B (accumulator[5]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (p_0[4]), .A (multiplicand[4]), .B (accumulator[4]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (p_0[3]), .A (multiplicand[3]), .B (accumulator[3]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (p_0[2]), .A (multiplicand[2]), .B (accumulator[2]), .CI (n_1));
FA_X1 i_1 (.CO (n_1), .S (p_0[1]), .A (multiplicand[1]), .B (accumulator[1]), .CI (n_0));
HA_X1 i_0 (.CO (n_0), .S (p_0[0]), .A (multiplicand[0]), .B (accumulator[0]));

endmodule //datapath__0_12

module datapath__0_10 (p_0, p_1);

output [63:0] p_0;
input [63:0] p_1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_65 (.ZN (n_33), .A (p_1[25]));
INV_X1 i_64 (.ZN (n_32), .A (p_1[21]));
INV_X1 i_63 (.ZN (n_31), .A (p_1[14]));
INV_X1 i_62 (.ZN (n_30), .A (p_1[11]));
OR3_X1 i_61 (.ZN (n_29), .A1 (p_1[2]), .A2 (p_1[1]), .A3 (p_1[0]));
OR2_X1 i_60 (.ZN (n_28), .A1 (n_29), .A2 (p_1[3]));
OR2_X1 i_59 (.ZN (n_27), .A1 (n_28), .A2 (p_1[4]));
OR3_X1 i_58 (.ZN (n_26), .A1 (n_27), .A2 (p_1[5]), .A3 (p_1[6]));
OR2_X1 i_57 (.ZN (n_25), .A1 (n_26), .A2 (p_1[7]));
OR3_X1 i_56 (.ZN (n_24), .A1 (n_25), .A2 (p_1[8]), .A3 (p_1[9]));
NOR2_X1 i_55 (.ZN (n_23), .A1 (n_24), .A2 (p_1[10]));
NAND2_X1 i_54 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_53 (.ZN (n_21), .A1 (n_22), .A2 (p_1[12]));
NOR3_X1 i_52 (.ZN (n_20), .A1 (n_22), .A2 (p_1[12]), .A3 (p_1[13]));
NAND2_X1 i_51 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_50 (.ZN (n_18), .A1 (n_19), .A2 (p_1[15]), .A3 (p_1[16]));
OR2_X1 i_49 (.ZN (n_17), .A1 (n_18), .A2 (p_1[17]));
NOR2_X1 i_48 (.ZN (n_16), .A1 (n_17), .A2 (p_1[18]));
NOR3_X1 i_47 (.ZN (n_15), .A1 (n_17), .A2 (p_1[18]), .A3 (p_1[19]));
NOR4_X1 i_46 (.ZN (n_14), .A1 (n_17), .A2 (p_1[18]), .A3 (p_1[19]), .A4 (p_1[20]));
NAND2_X1 i_45 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_44 (.ZN (n_12), .A1 (n_13), .A2 (p_1[22]));
NOR2_X1 i_43 (.ZN (n_11), .A1 (n_12), .A2 (p_1[23]));
NOR3_X1 i_42 (.ZN (n_10), .A1 (n_12), .A2 (p_1[23]), .A3 (p_1[24]));
NAND2_X1 i_41 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_40 (.ZN (n_8), .A1 (n_9), .A2 (p_1[26]), .A3 (p_1[27]));
NOR2_X1 i_39 (.ZN (n_7), .A1 (n_8), .A2 (p_1[28]));
NOR3_X1 i_38 (.ZN (n_6), .A1 (n_8), .A2 (p_1[28]), .A3 (p_1[29]));
NOR4_X2 i_37 (.ZN (n_5), .A1 (n_8), .A2 (p_1[28]), .A3 (p_1[29]), .A4 (p_1[30]));
NOR2_X4 i_36 (.ZN (p_0[63]), .A1 (p_1[31]), .A2 (n_5));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (p_1[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (p_1[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (p_1[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (p_1[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (p_1[27]), .B1 (n_9), .B2 (p_1[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (p_1[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (p_1[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (p_1[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (p_1[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (p_1[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (p_1[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (p_1[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (p_1[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (p_1[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (p_1[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (p_1[16]), .B1 (n_19), .B2 (p_1[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (p_1[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (p_1[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (p_1[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (p_1[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (p_1[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (p_1[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (p_1[9]), .B1 (n_25), .B2 (p_1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (p_1[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (p_1[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (p_1[6]), .B1 (n_27), .B2 (p_1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (p_1[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (p_1[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (p_1[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (p_1[2]), .B1 (p_1[1]), .B2 (p_1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (p_1[1]), .B (p_1[0]));

endmodule //datapath__0_10

module datapath (p_0, p_1);

output [31:0] p_0;
input [31:0] p_1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (p_1[25]));
INV_X1 i_63 (.ZN (n_32), .A (p_1[21]));
INV_X1 i_62 (.ZN (n_31), .A (p_1[14]));
INV_X1 i_61 (.ZN (n_30), .A (p_1[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (p_1[2]), .A2 (p_1[1]), .A3 (p_1[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (p_1[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (p_1[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (p_1[5]), .A3 (p_1[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (p_1[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (p_1[8]), .A3 (p_1[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (p_1[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (p_1[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (p_1[12]), .A3 (p_1[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (p_1[15]), .A3 (p_1[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (p_1[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (p_1[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (p_1[18]), .A3 (p_1[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (p_1[18]), .A3 (p_1[19]), .A4 (p_1[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (p_1[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (p_1[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (p_1[23]), .A3 (p_1[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (p_1[26]), .A3 (p_1[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (p_1[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (p_1[28]), .A3 (p_1[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (p_1[28]), .A3 (p_1[29]), .A4 (p_1[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (p_1[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (p_1[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (p_1[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (p_1[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (p_1[27]), .B1 (n_9), .B2 (p_1[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (p_1[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (p_1[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (p_1[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (p_1[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (p_1[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (p_1[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (p_1[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (p_1[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (p_1[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (p_1[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (p_1[16]), .B1 (n_19), .B2 (p_1[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (p_1[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (p_1[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (p_1[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (p_1[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (p_1[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (p_1[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (p_1[9]), .B1 (n_25), .B2 (p_1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (p_1[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (p_1[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (p_1[6]), .B1 (n_27), .B2 (p_1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (p_1[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (p_1[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (p_1[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (p_1[2]), .B1 (p_1[1]), .B2 (p_1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (p_1[1]), .B (p_1[0]));

endmodule //datapath

module sequential_multiplier (clk, rst, x, y, product);

output [63:0] product;
input clk;
input rst;
input [31:0] x;
input [31:0] y;
wire CTS_n_tid1_362;
wire CTS_n_tid0_299;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_0_104;
wire n_0_0_105;
wire n_0_0_0;
wire n_0_0_106;
wire n_0_0_1;
wire n_0_0_107;
wire n_0_0_2;
wire n_0_0_108;
wire n_0_0_109;
wire n_0_0_3;
wire n_0_368;
wire n_0_336;
wire n_0_337;
wire n_0_338;
wire n_0_339;
wire n_0_340;
wire n_0_341;
wire n_0_342;
wire n_0_343;
wire n_0_344;
wire n_0_345;
wire n_0_346;
wire n_0_347;
wire n_0_348;
wire n_0_349;
wire n_0_350;
wire n_0_351;
wire n_0_352;
wire n_0_353;
wire n_0_354;
wire n_0_355;
wire n_0_356;
wire n_0_357;
wire n_0_358;
wire n_0_359;
wire n_0_360;
wire n_0_361;
wire n_0_362;
wire n_0_363;
wire n_0_364;
wire n_0_365;
wire n_0_366;
wire n_0_367;
wire n_0_304;
wire n_0_305;
wire n_0_306;
wire n_0_307;
wire n_0_308;
wire n_0_309;
wire n_0_310;
wire n_0_311;
wire n_0_312;
wire n_0_313;
wire n_0_314;
wire n_0_315;
wire n_0_316;
wire n_0_317;
wire n_0_318;
wire n_0_319;
wire n_0_320;
wire n_0_321;
wire n_0_322;
wire n_0_323;
wire n_0_324;
wire n_0_325;
wire n_0_326;
wire n_0_327;
wire n_0_328;
wire n_0_329;
wire n_0_330;
wire n_0_331;
wire n_0_332;
wire n_0_333;
wire n_0_334;
wire n_0_335;
wire n_0_0_110;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_282;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_297;
wire n_0_298;
wire n_0_299;
wire n_0_300;
wire n_0_301;
wire n_0_302;
wire n_0_303;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_111;
wire n_0_0_112;
wire n_0_272;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_265;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_201;
wire n_0_0_37;
wire n_0_202;
wire n_0_0_38;
wire n_0_203;
wire n_0_0_39;
wire n_0_204;
wire n_0_0_40;
wire n_0_205;
wire n_0_0_41;
wire n_0_206;
wire n_0_0_42;
wire n_0_207;
wire n_0_0_43;
wire n_0_208;
wire n_0_0_44;
wire n_0_209;
wire n_0_0_45;
wire n_0_210;
wire n_0_0_46;
wire n_0_211;
wire n_0_0_47;
wire n_0_212;
wire n_0_0_48;
wire n_0_213;
wire n_0_0_49;
wire n_0_214;
wire n_0_0_50;
wire n_0_215;
wire n_0_0_51;
wire n_0_216;
wire n_0_0_52;
wire n_0_217;
wire n_0_0_53;
wire n_0_218;
wire n_0_0_54;
wire n_0_219;
wire n_0_0_55;
wire n_0_220;
wire n_0_0_56;
wire n_0_221;
wire n_0_0_57;
wire n_0_222;
wire n_0_0_58;
wire n_0_223;
wire n_0_0_59;
wire n_0_224;
wire n_0_0_60;
wire n_0_225;
wire n_0_0_61;
wire n_0_226;
wire n_0_0_62;
wire n_0_227;
wire n_0_0_63;
wire n_0_228;
wire n_0_0_64;
wire n_0_229;
wire n_0_0_65;
wire n_0_230;
wire n_0_0_66;
wire n_0_231;
wire n_0_0_67;
wire n_0_0_68;
wire n_0_232;
wire n_0_0_69;
wire n_0_233;
wire n_0_0_70;
wire n_0_234;
wire n_0_0_71;
wire n_0_235;
wire n_0_0_72;
wire n_0_236;
wire n_0_0_73;
wire n_0_237;
wire n_0_0_74;
wire n_0_238;
wire n_0_0_75;
wire n_0_239;
wire n_0_0_76;
wire n_0_240;
wire n_0_0_77;
wire n_0_241;
wire n_0_0_78;
wire n_0_242;
wire n_0_0_79;
wire n_0_243;
wire n_0_0_80;
wire n_0_244;
wire n_0_0_81;
wire n_0_245;
wire n_0_0_82;
wire n_0_246;
wire n_0_0_83;
wire n_0_247;
wire n_0_0_84;
wire n_0_248;
wire n_0_0_85;
wire n_0_249;
wire n_0_0_86;
wire n_0_250;
wire n_0_0_87;
wire n_0_251;
wire n_0_0_88;
wire n_0_252;
wire n_0_0_89;
wire n_0_253;
wire n_0_0_90;
wire n_0_254;
wire n_0_0_91;
wire n_0_255;
wire n_0_0_92;
wire n_0_256;
wire n_0_0_93;
wire n_0_257;
wire n_0_0_94;
wire n_0_258;
wire n_0_0_95;
wire n_0_259;
wire n_0_0_96;
wire n_0_260;
wire n_0_0_97;
wire n_0_261;
wire n_0_0_98;
wire n_0_262;
wire n_0_0_99;
wire n_0_263;
wire n_0_0_100;
wire n_0_264;
wire n_0_0_101;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_191;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_0_102;
wire n_0_0_113;
wire n_0_0_103;
wire n_0_369;
wire n_0_428;
wire n_0_429;
wire n_0_430;
wire n_0_431;
wire n_0_432;
wire n_0_433;
wire n_0_434;
wire n_0_435;
wire n_0_436;
wire n_0_437;
wire n_0_438;
wire n_0_439;
wire n_0_440;
wire n_0_441;
wire n_0_442;
wire n_0_443;
wire n_0_444;
wire n_0_445;
wire n_0_446;
wire n_0_447;
wire n_0_448;
wire n_0_449;
wire n_0_450;
wire n_0_451;
wire n_0_452;
wire n_0_453;
wire n_0_454;
wire n_0_455;
wire n_0_456;
wire n_0_457;
wire n_0_458;
wire n_0_459;
wire n_0_460;
wire n_0_461;
wire n_0_462;
wire n_0_463;
wire n_0_464;
wire n_0_465;
wire n_0_466;
wire n_0_467;
wire n_0_468;
wire n_0_469;
wire n_0_470;
wire n_0_471;
wire n_0_472;
wire n_0_473;
wire n_0_474;
wire n_0_475;
wire n_0_476;
wire n_0_477;
wire n_0_478;
wire n_0_479;
wire n_0_480;
wire n_0_481;
wire n_0_482;
wire n_0_483;
wire n_0_484;
wire n_0_485;
wire n_0_486;
wire n_0_487;
wire n_0_488;
wire n_0_489;
wire n_0_490;
wire n_0_372;
wire n_0_373;
wire n_0_374;
wire n_0_375;
wire n_0_376;
wire n_0_377;
wire n_0_378;
wire n_0_379;
wire n_0_380;
wire n_0_381;
wire n_0_382;
wire n_0_383;
wire n_0_384;
wire n_0_385;
wire n_0_386;
wire n_0_387;
wire n_0_388;
wire n_0_389;
wire n_0_390;
wire n_0_391;
wire n_0_392;
wire n_0_393;
wire n_0_394;
wire n_0_395;
wire n_0_396;
wire n_0_397;
wire n_0_398;
wire n_0_399;
wire n_0_400;
wire n_0_401;
wire n_0_402;
wire n_0_403;
wire n_0_404;
wire n_0_405;
wire n_0_406;
wire n_0_407;
wire n_0_408;
wire n_0_409;
wire n_0_410;
wire n_0_411;
wire n_0_412;
wire n_0_413;
wire n_0_414;
wire n_0_415;
wire n_0_416;
wire n_0_417;
wire n_0_418;
wire n_0_419;
wire n_0_420;
wire n_0_421;
wire n_0_422;
wire n_0_423;
wire n_0_424;
wire n_0_425;
wire n_0_426;
wire n_0_427;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire \ctr[5] ;
wire \ctr[4] ;
wire \ctr[3] ;
wire \ctr[2] ;
wire \ctr[1] ;
wire \ctr[0] ;
wire n_0_132;
wire \multiplier[31] ;
wire \multiplier[30] ;
wire \multiplier[29] ;
wire \multiplier[28] ;
wire \multiplier[27] ;
wire \multiplier[26] ;
wire \multiplier[25] ;
wire \multiplier[24] ;
wire \multiplier[23] ;
wire \multiplier[22] ;
wire \multiplier[21] ;
wire \multiplier[20] ;
wire \multiplier[19] ;
wire \multiplier[18] ;
wire \multiplier[17] ;
wire \multiplier[16] ;
wire \multiplier[15] ;
wire \multiplier[14] ;
wire \multiplier[13] ;
wire \multiplier[12] ;
wire \multiplier[11] ;
wire \multiplier[10] ;
wire \multiplier[9] ;
wire \multiplier[8] ;
wire \multiplier[7] ;
wire \multiplier[6] ;
wire \multiplier[5] ;
wire \multiplier[4] ;
wire \multiplier[3] ;
wire \multiplier[2] ;
wire \multiplier[1] ;
wire \multiplier[0] ;
wire uc_0;
wire uc_1;
wire uc_2;
wire uc_3;
wire uc_4;
wire uc_5;
wire uc_6;
wire uc_7;
wire uc_8;
wire uc_9;
wire uc_10;
wire uc_11;
wire uc_12;
wire uc_13;
wire uc_14;
wire uc_15;
wire uc_16;
wire uc_17;
wire uc_18;
wire uc_19;
wire uc_20;
wire uc_21;
wire uc_22;
wire uc_23;
wire uc_24;
wire uc_25;
wire uc_26;
wire uc_27;
wire uc_28;
wire uc_29;
wire uc_30;
wire uc_31;
wire uc_32;
wire uc_33;
wire uc_34;
wire uc_35;
wire uc_36;
wire uc_37;
wire uc_38;
wire uc_39;
wire uc_40;
wire uc_41;
wire uc_42;
wire uc_43;
wire uc_44;
wire uc_45;
wire uc_46;
wire uc_47;
wire uc_48;
wire uc_49;
wire uc_50;
wire uc_51;
wire uc_52;
wire uc_53;
wire uc_54;
wire uc_55;
wire uc_56;
wire uc_57;
wire uc_58;
wire uc_59;
wire uc_60;
wire uc_61;
wire uc_62;
wire uc_63;
wire uc_64;
wire hfn_ipo_n19;
wire hfn_ipo_n20;
wire hfn_ipo_n21;
wire hfn_ipo_n22;
wire hfn_ipo_n24;
wire hfn_ipo_n17;
wire hfn_ipo_n18;
wire drc_ipo_n25;
wire drc_ipo_n26;
wire drc_ipo_n27;
wire drc_ipo_n28;
wire drc_ipo_n29;
wire drc_ipo_n30;
wire drc_ipo_n31;
wire drc_ipo_n32;
wire drc_ipo_n33;
wire drc_ipo_n34;
wire drc_ipo_n35;
wire drc_ipo_n36;
wire drc_ipo_n37;
wire drc_ipo_n38;
wire drc_ipo_n39;
wire drc_ipo_n40;
wire drc_ipo_n41;
wire drc_ipo_n42;
wire drc_ipo_n43;
wire drc_ipo_n44;
wire drc_ipo_n45;
wire drc_ipo_n46;
wire drc_ipo_n47;
wire drc_ipo_n48;
wire drc_ipo_n49;
wire drc_ipo_n50;
wire drc_ipo_n51;
wire drc_ipo_n52;
wire drc_ipo_n53;
wire drc_ipo_n54;
wire drc_ipo_n55;
wire drc_ipo_n56;
wire drc_ipo_n57;
wire drc_ipo_n58;
wire drc_ipo_n59;
wire drc_ipo_n60;
wire drc_ipo_n61;
wire drc_ipo_n62;
wire drc_ipo_n63;
wire drc_ipo_n64;
wire drc_ipo_n65;
wire drc_ipo_n66;
wire drc_ipo_n67;
wire drc_ipo_n68;
wire drc_ipo_n69;
wire drc_ipo_n70;
wire drc_ipo_n71;
wire drc_ipo_n72;
wire drc_ipo_n73;
wire drc_ipo_n74;
wire drc_ipo_n75;
wire drc_ipo_n76;
wire drc_ipo_n77;
wire drc_ipo_n78;
wire drc_ipo_n79;
wire drc_ipo_n80;
wire drc_ipo_n81;
wire drc_ipo_n82;
wire drc_ipo_n83;
wire drc_ipo_n84;
wire drc_ipo_n85;
wire drc_ipo_n86;
wire drc_ipo_n87;
wire drc_ipo_n88;
wire drc_ipo_n89;
wire CTS_n_tid0_300;
wire CTS_n_tid1_126;
wire CTS_n_tid0_128;
wire CTS_n_tid0_129;
wire CTS_n_tid1_130;
wire CTS_n_tid0_132;
wire CTS_n_tid0_133;
wire CTS_n_tid0_285;


CLKGATETST_X4 clk_gate_multiplicand_reg (.GCK (CTS_n_tid0_285), .CK (CTS_n_tid1_362)
    , .E (n_0_265), .SE (1'b0 ));
DFF_X1 \multiplier_reg[0]  (.Q (\multiplier[0] ), .CK (n_0_132), .D (n_0_336));
DFF_X1 \multiplier_reg[1]  (.Q (\multiplier[1] ), .CK (n_0_132), .D (n_0_273));
DFF_X1 \multiplier_reg[2]  (.Q (\multiplier[2] ), .CK (n_0_132), .D (n_0_274));
DFF_X1 \multiplier_reg[3]  (.Q (\multiplier[3] ), .CK (n_0_132), .D (n_0_275));
DFF_X1 \multiplier_reg[4]  (.Q (\multiplier[4] ), .CK (n_0_132), .D (n_0_276));
DFF_X1 \multiplier_reg[5]  (.Q (\multiplier[5] ), .CK (n_0_132), .D (n_0_277));
DFF_X1 \multiplier_reg[6]  (.Q (\multiplier[6] ), .CK (n_0_132), .D (n_0_278));
DFF_X1 \multiplier_reg[7]  (.Q (\multiplier[7] ), .CK (n_0_132), .D (n_0_279));
DFF_X1 \multiplier_reg[8]  (.Q (\multiplier[8] ), .CK (n_0_132), .D (n_0_280));
DFF_X1 \multiplier_reg[9]  (.Q (\multiplier[9] ), .CK (n_0_132), .D (n_0_281));
DFF_X1 \multiplier_reg[10]  (.Q (\multiplier[10] ), .CK (n_0_132), .D (n_0_282));
DFF_X1 \multiplier_reg[11]  (.Q (\multiplier[11] ), .CK (n_0_132), .D (n_0_283));
DFF_X1 \multiplier_reg[12]  (.Q (\multiplier[12] ), .CK (n_0_132), .D (n_0_284));
DFF_X1 \multiplier_reg[13]  (.Q (\multiplier[13] ), .CK (n_0_132), .D (n_0_285));
DFF_X1 \multiplier_reg[14]  (.Q (\multiplier[14] ), .CK (n_0_132), .D (n_0_286));
DFF_X1 \multiplier_reg[15]  (.Q (\multiplier[15] ), .CK (n_0_132), .D (n_0_287));
DFF_X1 \multiplier_reg[16]  (.Q (\multiplier[16] ), .CK (n_0_132), .D (n_0_288));
DFF_X1 \multiplier_reg[17]  (.Q (\multiplier[17] ), .CK (n_0_132), .D (n_0_289));
DFF_X1 \multiplier_reg[18]  (.Q (\multiplier[18] ), .CK (n_0_132), .D (n_0_290));
DFF_X1 \multiplier_reg[19]  (.Q (\multiplier[19] ), .CK (n_0_132), .D (n_0_291));
DFF_X1 \multiplier_reg[20]  (.Q (\multiplier[20] ), .CK (n_0_132), .D (n_0_292));
DFF_X1 \multiplier_reg[21]  (.Q (\multiplier[21] ), .CK (n_0_132), .D (n_0_293));
DFF_X1 \multiplier_reg[22]  (.Q (\multiplier[22] ), .CK (n_0_132), .D (n_0_294));
DFF_X1 \multiplier_reg[23]  (.Q (\multiplier[23] ), .CK (n_0_132), .D (n_0_295));
DFF_X1 \multiplier_reg[24]  (.Q (\multiplier[24] ), .CK (n_0_132), .D (n_0_296));
DFF_X1 \multiplier_reg[25]  (.Q (\multiplier[25] ), .CK (n_0_132), .D (n_0_297));
DFF_X1 \multiplier_reg[26]  (.Q (\multiplier[26] ), .CK (n_0_132), .D (n_0_298));
DFF_X1 \multiplier_reg[27]  (.Q (\multiplier[27] ), .CK (n_0_132), .D (n_0_299));
DFF_X1 \multiplier_reg[28]  (.Q (\multiplier[28] ), .CK (n_0_132), .D (n_0_300));
DFF_X1 \multiplier_reg[29]  (.Q (\multiplier[29] ), .CK (n_0_132), .D (n_0_301));
DFF_X1 \multiplier_reg[30]  (.Q (\multiplier[30] ), .CK (n_0_132), .D (n_0_302));
DFF_X1 \multiplier_reg[31]  (.Q (\multiplier[31] ), .CK (n_0_132), .D (n_0_303));
CLKGATETST_X1 clk_gate_multiplier_reg (.GCK (n_0_132), .CK (CTS_n_tid1_362), .E (drc_ipo_n89), .SE (1'b0 ));
DFF_X1 \ctr_reg[0]  (.Q (\ctr[0] ), .CK (CTS_n_tid0_129), .D (n_0_266));
DFF_X1 \ctr_reg[1]  (.Q (\ctr[1] ), .CK (CTS_n_tid0_129), .D (n_0_267));
DFF_X1 \ctr_reg[2]  (.Q (\ctr[2] ), .CK (CTS_n_tid0_129), .D (n_0_268));
DFF_X1 \ctr_reg[3]  (.Q (\ctr[3] ), .CK (CTS_n_tid0_129), .D (n_0_269));
DFF_X1 \ctr_reg[4]  (.Q (\ctr[4] ), .CK (CTS_n_tid0_129), .D (n_0_270));
DFF_X1 \ctr_reg[5]  (.Q (\ctr[5] ), .CK (CTS_n_tid0_129), .D (n_0_271));
DFF_X1 \accumulator_reg[0]  (.Q (n_0_8), .CK (CTS_n_tid1_126), .D (n_0_137));
DFF_X1 \accumulator_reg[1]  (.Q (n_0_7), .CK (CTS_n_tid1_126), .D (n_0_138));
DFF_X1 \accumulator_reg[2]  (.Q (n_0_6), .CK (CTS_n_tid1_126), .D (n_0_139));
DFF_X1 \accumulator_reg[3]  (.Q (n_0_5), .CK (CTS_n_tid1_126), .D (n_0_140));
DFF_X1 \accumulator_reg[4]  (.Q (n_0_4), .CK (CTS_n_tid1_126), .D (n_0_141));
DFF_X1 \accumulator_reg[5]  (.Q (n_0_3), .CK (CTS_n_tid1_126), .D (n_0_142));
DFF_X1 \accumulator_reg[6]  (.Q (n_0_2), .CK (CTS_n_tid1_126), .D (n_0_143));
DFF_X1 \accumulator_reg[7]  (.Q (n_0_1), .CK (CTS_n_tid1_126), .D (n_0_144));
DFF_X1 \accumulator_reg[8]  (.Q (n_0_427), .CK (CTS_n_tid1_126), .D (n_0_145));
DFF_X1 \accumulator_reg[9]  (.Q (n_0_426), .CK (CTS_n_tid1_126), .D (n_0_146));
DFF_X1 \accumulator_reg[10]  (.Q (n_0_425), .CK (CTS_n_tid1_126), .D (n_0_147));
DFF_X1 \accumulator_reg[11]  (.Q (n_0_424), .CK (CTS_n_tid1_126), .D (n_0_148));
DFF_X1 \accumulator_reg[12]  (.Q (n_0_423), .CK (CTS_n_tid1_126), .D (n_0_149));
DFF_X1 \accumulator_reg[13]  (.Q (n_0_422), .CK (CTS_n_tid1_126), .D (n_0_150));
DFF_X1 \accumulator_reg[14]  (.Q (n_0_421), .CK (CTS_n_tid1_126), .D (n_0_151));
DFF_X1 \accumulator_reg[15]  (.Q (n_0_420), .CK (CTS_n_tid1_126), .D (n_0_152));
DFF_X1 \accumulator_reg[16]  (.Q (n_0_419), .CK (CTS_n_tid1_126), .D (n_0_153));
DFF_X1 \accumulator_reg[17]  (.Q (n_0_418), .CK (CTS_n_tid1_126), .D (n_0_154));
DFF_X1 \accumulator_reg[18]  (.Q (n_0_417), .CK (CTS_n_tid1_126), .D (n_0_155));
DFF_X1 \accumulator_reg[19]  (.Q (n_0_416), .CK (CTS_n_tid1_126), .D (n_0_156));
DFF_X1 \accumulator_reg[20]  (.Q (n_0_415), .CK (CTS_n_tid1_126), .D (n_0_157));
DFF_X1 \accumulator_reg[21]  (.Q (n_0_414), .CK (CTS_n_tid1_126), .D (n_0_158));
DFF_X1 \accumulator_reg[22]  (.Q (n_0_413), .CK (CTS_n_tid1_126), .D (n_0_159));
DFF_X1 \accumulator_reg[23]  (.Q (n_0_412), .CK (CTS_n_tid1_126), .D (n_0_160));
DFF_X1 \accumulator_reg[24]  (.Q (n_0_411), .CK (CTS_n_tid1_126), .D (n_0_161));
DFF_X1 \accumulator_reg[25]  (.Q (n_0_410), .CK (CTS_n_tid1_126), .D (n_0_162));
DFF_X1 \accumulator_reg[26]  (.Q (n_0_409), .CK (CTS_n_tid1_126), .D (n_0_163));
DFF_X1 \accumulator_reg[27]  (.Q (n_0_408), .CK (CTS_n_tid1_126), .D (n_0_164));
DFF_X1 \accumulator_reg[28]  (.Q (n_0_407), .CK (CTS_n_tid1_126), .D (n_0_165));
DFF_X1 \accumulator_reg[29]  (.Q (n_0_406), .CK (CTS_n_tid1_126), .D (n_0_166));
DFF_X1 \accumulator_reg[30]  (.Q (n_0_405), .CK (CTS_n_tid1_126), .D (n_0_167));
DFF_X1 \accumulator_reg[31]  (.Q (n_0_404), .CK (CTS_n_tid1_126), .D (n_0_168));
DFF_X1 \accumulator_reg[32]  (.Q (n_0_403), .CK (CTS_n_tid1_126), .D (n_0_169));
DFF_X1 \accumulator_reg[33]  (.Q (n_0_402), .CK (CTS_n_tid1_126), .D (n_0_170));
DFF_X1 \accumulator_reg[34]  (.Q (n_0_401), .CK (CTS_n_tid1_126), .D (n_0_171));
DFF_X1 \accumulator_reg[35]  (.Q (n_0_400), .CK (CTS_n_tid1_126), .D (n_0_172));
DFF_X1 \accumulator_reg[36]  (.Q (n_0_399), .CK (CTS_n_tid1_126), .D (n_0_173));
DFF_X1 \accumulator_reg[37]  (.Q (n_0_398), .CK (CTS_n_tid1_126), .D (n_0_174));
DFF_X1 \accumulator_reg[38]  (.Q (n_0_397), .CK (CTS_n_tid1_126), .D (n_0_175));
DFF_X1 \accumulator_reg[39]  (.Q (n_0_396), .CK (CTS_n_tid1_126), .D (n_0_176));
DFF_X1 \accumulator_reg[40]  (.Q (n_0_395), .CK (CTS_n_tid1_126), .D (n_0_177));
DFF_X1 \accumulator_reg[41]  (.Q (n_0_394), .CK (CTS_n_tid1_126), .D (n_0_178));
DFF_X1 \accumulator_reg[42]  (.Q (n_0_393), .CK (CTS_n_tid1_126), .D (n_0_179));
DFF_X1 \accumulator_reg[43]  (.Q (n_0_392), .CK (CTS_n_tid1_126), .D (n_0_180));
DFF_X1 \accumulator_reg[44]  (.Q (n_0_391), .CK (CTS_n_tid1_126), .D (n_0_181));
DFF_X1 \accumulator_reg[45]  (.Q (n_0_390), .CK (CTS_n_tid1_126), .D (n_0_182));
DFF_X1 \accumulator_reg[46]  (.Q (n_0_389), .CK (CTS_n_tid1_126), .D (n_0_183));
DFF_X1 \accumulator_reg[47]  (.Q (n_0_388), .CK (CTS_n_tid1_126), .D (n_0_184));
DFF_X1 \accumulator_reg[48]  (.Q (n_0_387), .CK (CTS_n_tid1_126), .D (n_0_185));
DFF_X1 \accumulator_reg[49]  (.Q (n_0_386), .CK (CTS_n_tid1_126), .D (n_0_186));
DFF_X1 \accumulator_reg[50]  (.Q (n_0_385), .CK (CTS_n_tid1_126), .D (n_0_187));
DFF_X1 \accumulator_reg[51]  (.Q (n_0_384), .CK (CTS_n_tid1_126), .D (n_0_188));
DFF_X1 \accumulator_reg[52]  (.Q (n_0_383), .CK (CTS_n_tid1_126), .D (n_0_189));
DFF_X1 \accumulator_reg[53]  (.Q (n_0_382), .CK (CTS_n_tid1_126), .D (n_0_190));
DFF_X1 \accumulator_reg[54]  (.Q (n_0_381), .CK (CTS_n_tid1_126), .D (n_0_191));
DFF_X1 \accumulator_reg[55]  (.Q (n_0_380), .CK (CTS_n_tid1_126), .D (n_0_192));
DFF_X1 \accumulator_reg[56]  (.Q (n_0_379), .CK (CTS_n_tid1_126), .D (n_0_193));
DFF_X1 \accumulator_reg[57]  (.Q (n_0_378), .CK (CTS_n_tid1_126), .D (n_0_194));
DFF_X1 \accumulator_reg[58]  (.Q (n_0_377), .CK (CTS_n_tid1_126), .D (n_0_195));
DFF_X1 \accumulator_reg[59]  (.Q (n_0_376), .CK (CTS_n_tid1_126), .D (n_0_196));
DFF_X1 \accumulator_reg[60]  (.Q (n_0_375), .CK (CTS_n_tid1_126), .D (n_0_197));
DFF_X1 \accumulator_reg[61]  (.Q (n_0_374), .CK (CTS_n_tid1_126), .D (n_0_198));
DFF_X1 \accumulator_reg[62]  (.Q (n_0_373), .CK (CTS_n_tid1_126), .D (n_0_199));
DFF_X1 \accumulator_reg[63]  (.Q (n_0_372), .CK (CTS_n_tid1_126), .D (n_0_200));
CLKGATETST_X8 clk_gate_accumulator_reg (.GCK (CTS_n_tid1_130), .CK (CTS_n_tid1_362)
    , .E (n_0_272), .SE (1'b0 ));
DFF_X1 \multiplicand_reg[0]  (.Q (n_0_490), .CK (CTS_n_tid0_129), .D (n_0_201));
DFF_X1 \multiplicand_reg[1]  (.Q (n_0_489), .CK (CTS_n_tid0_129), .D (n_0_202));
DFF_X1 \multiplicand_reg[2]  (.Q (n_0_488), .CK (CTS_n_tid0_129), .D (n_0_203));
DFF_X1 \multiplicand_reg[3]  (.Q (n_0_487), .CK (CTS_n_tid0_132), .D (n_0_204));
DFF_X1 \multiplicand_reg[4]  (.Q (n_0_486), .CK (CTS_n_tid0_132), .D (n_0_205));
DFF_X1 \multiplicand_reg[5]  (.Q (n_0_485), .CK (CTS_n_tid0_132), .D (n_0_206));
DFF_X1 \multiplicand_reg[6]  (.Q (n_0_484), .CK (CTS_n_tid0_132), .D (n_0_207));
DFF_X1 \multiplicand_reg[7]  (.Q (n_0_483), .CK (CTS_n_tid0_132), .D (n_0_208));
DFF_X1 \multiplicand_reg[8]  (.Q (n_0_482), .CK (CTS_n_tid0_132), .D (n_0_209));
DFF_X1 \multiplicand_reg[9]  (.Q (n_0_481), .CK (CTS_n_tid0_132), .D (n_0_210));
DFF_X1 \multiplicand_reg[10]  (.Q (n_0_480), .CK (CTS_n_tid0_132), .D (n_0_211));
DFF_X1 \multiplicand_reg[11]  (.Q (n_0_479), .CK (CTS_n_tid0_133), .D (n_0_212));
DFF_X1 \multiplicand_reg[12]  (.Q (n_0_478), .CK (CTS_n_tid0_133), .D (n_0_213));
DFF_X1 \multiplicand_reg[13]  (.Q (n_0_477), .CK (CTS_n_tid0_133), .D (n_0_214));
DFF_X1 \multiplicand_reg[14]  (.Q (n_0_476), .CK (CTS_n_tid0_133), .D (n_0_215));
DFF_X1 \multiplicand_reg[15]  (.Q (n_0_475), .CK (CTS_n_tid0_133), .D (n_0_216));
DFF_X1 \multiplicand_reg[16]  (.Q (n_0_474), .CK (CTS_n_tid0_133), .D (n_0_217));
DFF_X1 \multiplicand_reg[17]  (.Q (n_0_473), .CK (CTS_n_tid0_133), .D (n_0_218));
DFF_X1 \multiplicand_reg[18]  (.Q (n_0_472), .CK (CTS_n_tid0_133), .D (n_0_219));
DFF_X1 \multiplicand_reg[19]  (.Q (n_0_471), .CK (CTS_n_tid0_133), .D (n_0_220));
DFF_X1 \multiplicand_reg[20]  (.Q (n_0_470), .CK (CTS_n_tid0_133), .D (n_0_221));
DFF_X1 \multiplicand_reg[21]  (.Q (n_0_469), .CK (CTS_n_tid0_133), .D (n_0_222));
DFF_X1 \multiplicand_reg[22]  (.Q (n_0_468), .CK (CTS_n_tid0_133), .D (n_0_223));
DFF_X1 \multiplicand_reg[23]  (.Q (n_0_467), .CK (CTS_n_tid0_133), .D (n_0_224));
DFF_X1 \multiplicand_reg[24]  (.Q (n_0_466), .CK (CTS_n_tid0_133), .D (n_0_225));
DFF_X1 \multiplicand_reg[25]  (.Q (n_0_465), .CK (CTS_n_tid0_133), .D (n_0_226));
DFF_X1 \multiplicand_reg[26]  (.Q (n_0_464), .CK (CTS_n_tid0_133), .D (n_0_227));
DFF_X1 \multiplicand_reg[27]  (.Q (n_0_463), .CK (CTS_n_tid0_133), .D (n_0_228));
DFF_X1 \multiplicand_reg[28]  (.Q (n_0_462), .CK (CTS_n_tid0_133), .D (n_0_229));
DFF_X1 \multiplicand_reg[29]  (.Q (n_0_461), .CK (CTS_n_tid0_133), .D (n_0_230));
DFF_X1 \multiplicand_reg[30]  (.Q (n_0_460), .CK (CTS_n_tid0_133), .D (n_0_231));
DFF_X1 \multiplicand_reg[31]  (.Q (n_0_459), .CK (CTS_n_tid0_132), .D (n_0_232));
DFF_X1 \multiplicand_reg[32]  (.Q (n_0_458), .CK (CTS_n_tid0_132), .D (n_0_233));
DFF_X1 \multiplicand_reg[33]  (.Q (n_0_457), .CK (CTS_n_tid0_132), .D (n_0_234));
DFF_X1 \multiplicand_reg[34]  (.Q (n_0_456), .CK (CTS_n_tid0_132), .D (n_0_235));
DFF_X1 \multiplicand_reg[35]  (.Q (n_0_455), .CK (CTS_n_tid0_128), .D (n_0_236));
DFF_X1 \multiplicand_reg[36]  (.Q (n_0_454), .CK (CTS_n_tid0_128), .D (n_0_237));
DFF_X1 \multiplicand_reg[37]  (.Q (n_0_453), .CK (CTS_n_tid0_128), .D (n_0_238));
DFF_X1 \multiplicand_reg[38]  (.Q (n_0_452), .CK (CTS_n_tid0_128), .D (n_0_239));
DFF_X1 \multiplicand_reg[39]  (.Q (n_0_451), .CK (CTS_n_tid0_128), .D (n_0_240));
DFF_X1 \multiplicand_reg[40]  (.Q (n_0_450), .CK (CTS_n_tid0_128), .D (n_0_241));
DFF_X1 \multiplicand_reg[41]  (.Q (n_0_449), .CK (CTS_n_tid0_132), .D (n_0_242));
DFF_X1 \multiplicand_reg[42]  (.Q (n_0_448), .CK (CTS_n_tid0_132), .D (n_0_243));
DFF_X1 \multiplicand_reg[43]  (.Q (n_0_447), .CK (CTS_n_tid0_132), .D (n_0_244));
DFF_X1 \multiplicand_reg[44]  (.Q (n_0_446), .CK (CTS_n_tid0_132), .D (n_0_245));
DFF_X1 \multiplicand_reg[45]  (.Q (n_0_445), .CK (CTS_n_tid0_132), .D (n_0_246));
DFF_X1 \multiplicand_reg[46]  (.Q (n_0_444), .CK (CTS_n_tid0_132), .D (n_0_247));
DFF_X1 \multiplicand_reg[47]  (.Q (n_0_443), .CK (CTS_n_tid0_132), .D (n_0_248));
DFF_X1 \multiplicand_reg[48]  (.Q (n_0_442), .CK (CTS_n_tid0_128), .D (n_0_249));
DFF_X1 \multiplicand_reg[49]  (.Q (n_0_441), .CK (CTS_n_tid0_128), .D (n_0_250));
DFF_X1 \multiplicand_reg[50]  (.Q (n_0_440), .CK (CTS_n_tid0_128), .D (n_0_251));
DFF_X1 \multiplicand_reg[51]  (.Q (n_0_439), .CK (CTS_n_tid0_128), .D (n_0_252));
DFF_X1 \multiplicand_reg[52]  (.Q (n_0_438), .CK (CTS_n_tid0_128), .D (n_0_253));
DFF_X1 \multiplicand_reg[53]  (.Q (n_0_437), .CK (CTS_n_tid0_128), .D (n_0_254));
DFF_X1 \multiplicand_reg[54]  (.Q (n_0_436), .CK (CTS_n_tid0_128), .D (n_0_255));
DFF_X1 \multiplicand_reg[55]  (.Q (n_0_435), .CK (CTS_n_tid0_128), .D (n_0_256));
DFF_X1 \multiplicand_reg[56]  (.Q (n_0_434), .CK (CTS_n_tid0_128), .D (n_0_257));
DFF_X1 \multiplicand_reg[57]  (.Q (n_0_433), .CK (CTS_n_tid0_128), .D (n_0_258));
DFF_X1 \multiplicand_reg[58]  (.Q (n_0_432), .CK (CTS_n_tid0_128), .D (n_0_259));
DFF_X1 \multiplicand_reg[59]  (.Q (n_0_431), .CK (CTS_n_tid0_129), .D (n_0_260));
DFF_X1 \multiplicand_reg[60]  (.Q (n_0_430), .CK (CTS_n_tid0_129), .D (n_0_261));
DFF_X1 \multiplicand_reg[61]  (.Q (n_0_429), .CK (CTS_n_tid0_129), .D (n_0_262));
DFF_X1 \multiplicand_reg[62]  (.Q (n_0_428), .CK (CTS_n_tid0_129), .D (n_0_263));
DFF_X1 \multiplicand_reg[63]  (.Q (n_0_369), .CK (CTS_n_tid0_129), .D (n_0_264));
INV_X1 i_0_0_341 (.ZN (n_0_0_103), .A (drc_ipo_n89));
INV_X2 i_0_0_340 (.ZN (n_0_0_113), .A (hfn_ipo_n20));
INV_X1 i_0_0_339 (.ZN (n_0_0_102), .A (\ctr[5] ));
AND2_X1 i_0_0_338 (.ZN (n_0_200), .A1 (n_0_0_103), .A2 (n_0_136));
AND2_X1 i_0_0_337 (.ZN (n_0_199), .A1 (n_0_0_103), .A2 (n_0_135));
AND2_X1 i_0_0_336 (.ZN (n_0_198), .A1 (n_0_0_103), .A2 (n_0_134));
AND2_X1 i_0_0_335 (.ZN (n_0_197), .A1 (n_0_0_103), .A2 (n_0_133));
AND2_X1 i_0_0_334 (.ZN (n_0_196), .A1 (n_0_0_103), .A2 (n_0_131));
AND2_X1 i_0_0_333 (.ZN (n_0_195), .A1 (n_0_0_103), .A2 (n_0_130));
AND2_X1 i_0_0_332 (.ZN (n_0_194), .A1 (n_0_0_103), .A2 (n_0_129));
AND2_X1 i_0_0_331 (.ZN (n_0_193), .A1 (n_0_0_103), .A2 (n_0_128));
AND2_X1 i_0_0_330 (.ZN (n_0_192), .A1 (n_0_0_103), .A2 (n_0_127));
AND2_X1 i_0_0_329 (.ZN (n_0_191), .A1 (n_0_0_103), .A2 (n_0_126));
AND2_X1 i_0_0_328 (.ZN (n_0_190), .A1 (n_0_0_103), .A2 (n_0_125));
AND2_X1 i_0_0_327 (.ZN (n_0_189), .A1 (n_0_0_103), .A2 (n_0_124));
AND2_X1 i_0_0_326 (.ZN (n_0_188), .A1 (n_0_0_103), .A2 (n_0_123));
AND2_X1 i_0_0_325 (.ZN (n_0_187), .A1 (n_0_0_103), .A2 (n_0_122));
AND2_X1 i_0_0_324 (.ZN (n_0_186), .A1 (n_0_0_103), .A2 (n_0_121));
AND2_X1 i_0_0_323 (.ZN (n_0_185), .A1 (n_0_0_103), .A2 (n_0_120));
AND2_X1 i_0_0_322 (.ZN (n_0_184), .A1 (hfn_ipo_n24), .A2 (n_0_119));
AND2_X1 i_0_0_321 (.ZN (n_0_183), .A1 (hfn_ipo_n24), .A2 (n_0_118));
AND2_X1 i_0_0_320 (.ZN (n_0_182), .A1 (hfn_ipo_n24), .A2 (n_0_117));
AND2_X1 i_0_0_319 (.ZN (n_0_181), .A1 (hfn_ipo_n24), .A2 (n_0_116));
AND2_X1 i_0_0_318 (.ZN (n_0_180), .A1 (hfn_ipo_n24), .A2 (n_0_115));
AND2_X1 i_0_0_317 (.ZN (n_0_179), .A1 (hfn_ipo_n24), .A2 (n_0_114));
AND2_X1 i_0_0_316 (.ZN (n_0_178), .A1 (hfn_ipo_n24), .A2 (n_0_113));
AND2_X1 i_0_0_315 (.ZN (n_0_177), .A1 (hfn_ipo_n24), .A2 (n_0_112));
AND2_X1 i_0_0_314 (.ZN (n_0_176), .A1 (n_0_0_103), .A2 (n_0_111));
AND2_X1 i_0_0_313 (.ZN (n_0_175), .A1 (n_0_0_103), .A2 (n_0_110));
AND2_X1 i_0_0_312 (.ZN (n_0_174), .A1 (n_0_0_103), .A2 (n_0_109));
AND2_X1 i_0_0_311 (.ZN (n_0_173), .A1 (n_0_0_103), .A2 (n_0_108));
AND2_X1 i_0_0_310 (.ZN (n_0_172), .A1 (n_0_0_103), .A2 (n_0_107));
AND2_X1 i_0_0_309 (.ZN (n_0_171), .A1 (hfn_ipo_n24), .A2 (n_0_106));
AND2_X1 i_0_0_308 (.ZN (n_0_170), .A1 (hfn_ipo_n24), .A2 (n_0_105));
AND2_X1 i_0_0_307 (.ZN (n_0_169), .A1 (hfn_ipo_n24), .A2 (n_0_104));
AND2_X1 i_0_0_306 (.ZN (n_0_168), .A1 (hfn_ipo_n24), .A2 (n_0_103));
AND2_X1 i_0_0_305 (.ZN (n_0_167), .A1 (hfn_ipo_n24), .A2 (n_0_102));
AND2_X1 i_0_0_304 (.ZN (n_0_166), .A1 (hfn_ipo_n24), .A2 (n_0_101));
AND2_X1 i_0_0_303 (.ZN (n_0_165), .A1 (hfn_ipo_n24), .A2 (n_0_100));
AND2_X1 i_0_0_302 (.ZN (n_0_164), .A1 (hfn_ipo_n24), .A2 (n_0_99));
AND2_X1 i_0_0_301 (.ZN (n_0_163), .A1 (hfn_ipo_n24), .A2 (n_0_98));
AND2_X1 i_0_0_300 (.ZN (n_0_162), .A1 (hfn_ipo_n24), .A2 (n_0_97));
AND2_X1 i_0_0_299 (.ZN (n_0_161), .A1 (hfn_ipo_n24), .A2 (n_0_96));
AND2_X1 i_0_0_298 (.ZN (n_0_160), .A1 (hfn_ipo_n24), .A2 (n_0_95));
AND2_X1 i_0_0_297 (.ZN (n_0_159), .A1 (hfn_ipo_n24), .A2 (n_0_94));
AND2_X1 i_0_0_296 (.ZN (n_0_158), .A1 (hfn_ipo_n24), .A2 (n_0_93));
AND2_X1 i_0_0_295 (.ZN (n_0_157), .A1 (hfn_ipo_n24), .A2 (n_0_92));
AND2_X1 i_0_0_294 (.ZN (n_0_156), .A1 (hfn_ipo_n24), .A2 (n_0_91));
AND2_X1 i_0_0_293 (.ZN (n_0_155), .A1 (hfn_ipo_n24), .A2 (n_0_90));
AND2_X1 i_0_0_292 (.ZN (n_0_154), .A1 (hfn_ipo_n24), .A2 (n_0_89));
AND2_X1 i_0_0_291 (.ZN (n_0_153), .A1 (hfn_ipo_n24), .A2 (n_0_88));
AND2_X1 i_0_0_290 (.ZN (n_0_152), .A1 (hfn_ipo_n24), .A2 (n_0_87));
AND2_X1 i_0_0_289 (.ZN (n_0_151), .A1 (hfn_ipo_n24), .A2 (n_0_86));
AND2_X1 i_0_0_288 (.ZN (n_0_150), .A1 (hfn_ipo_n24), .A2 (n_0_85));
AND2_X1 i_0_0_287 (.ZN (n_0_149), .A1 (hfn_ipo_n24), .A2 (n_0_84));
AND2_X1 i_0_0_286 (.ZN (n_0_148), .A1 (hfn_ipo_n24), .A2 (n_0_83));
AND2_X1 i_0_0_285 (.ZN (n_0_147), .A1 (hfn_ipo_n24), .A2 (n_0_82));
AND2_X1 i_0_0_284 (.ZN (n_0_146), .A1 (hfn_ipo_n24), .A2 (n_0_81));
AND2_X1 i_0_0_283 (.ZN (n_0_145), .A1 (hfn_ipo_n24), .A2 (n_0_80));
AND2_X1 i_0_0_282 (.ZN (n_0_144), .A1 (hfn_ipo_n24), .A2 (n_0_79));
AND2_X1 i_0_0_281 (.ZN (n_0_143), .A1 (hfn_ipo_n24), .A2 (n_0_78));
AND2_X1 i_0_0_280 (.ZN (n_0_142), .A1 (hfn_ipo_n24), .A2 (n_0_77));
AND2_X1 i_0_0_279 (.ZN (n_0_141), .A1 (hfn_ipo_n24), .A2 (n_0_76));
AND2_X1 i_0_0_278 (.ZN (n_0_140), .A1 (hfn_ipo_n24), .A2 (n_0_75));
AND2_X1 i_0_0_277 (.ZN (n_0_139), .A1 (hfn_ipo_n24), .A2 (n_0_74));
AND2_X1 i_0_0_276 (.ZN (n_0_138), .A1 (hfn_ipo_n24), .A2 (n_0_73));
AND2_X1 i_0_0_275 (.ZN (n_0_137), .A1 (n_0_0_103), .A2 (n_0_72));
OAI21_X1 i_0_0_274 (.ZN (n_0_0_101), .A (n_0_304), .B1 (n_0_0_35), .B2 (hfn_ipo_n20));
INV_X1 i_0_0_273 (.ZN (n_0_264), .A (n_0_0_100));
AOI221_X1 i_0_0_272 (.ZN (n_0_0_100), .A (n_0_0_67), .B1 (hfn_ipo_n22), .B2 (n_0_428)
    , .C1 (hfn_ipo_n20), .C2 (n_0_71));
INV_X1 i_0_0_271 (.ZN (n_0_263), .A (n_0_0_99));
AOI221_X1 i_0_0_270 (.ZN (n_0_0_99), .A (n_0_0_67), .B1 (hfn_ipo_n22), .B2 (n_0_429)
    , .C1 (hfn_ipo_n20), .C2 (n_0_71));
INV_X1 i_0_0_269 (.ZN (n_0_262), .A (n_0_0_98));
AOI221_X1 i_0_0_268 (.ZN (n_0_0_98), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_430)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_267 (.ZN (n_0_261), .A (n_0_0_97));
AOI221_X1 i_0_0_266 (.ZN (n_0_0_97), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_431)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_265 (.ZN (n_0_260), .A (n_0_0_96));
AOI221_X1 i_0_0_264 (.ZN (n_0_0_96), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_432)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_263 (.ZN (n_0_259), .A (n_0_0_95));
AOI221_X1 i_0_0_262 (.ZN (n_0_0_95), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_433)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_261 (.ZN (n_0_258), .A (n_0_0_94));
AOI221_X1 i_0_0_260 (.ZN (n_0_0_94), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_434)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_259 (.ZN (n_0_257), .A (n_0_0_93));
AOI221_X1 i_0_0_258 (.ZN (n_0_0_93), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_435)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_257 (.ZN (n_0_256), .A (n_0_0_92));
AOI221_X1 i_0_0_256 (.ZN (n_0_0_92), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_436)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_255 (.ZN (n_0_255), .A (n_0_0_91));
AOI221_X1 i_0_0_254 (.ZN (n_0_0_91), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_437)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_253 (.ZN (n_0_254), .A (n_0_0_90));
AOI221_X1 i_0_0_252 (.ZN (n_0_0_90), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_438)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_251 (.ZN (n_0_253), .A (n_0_0_89));
AOI221_X1 i_0_0_250 (.ZN (n_0_0_89), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_439)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_249 (.ZN (n_0_252), .A (n_0_0_88));
AOI221_X1 i_0_0_248 (.ZN (n_0_0_88), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_440)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_247 (.ZN (n_0_251), .A (n_0_0_87));
AOI221_X1 i_0_0_246 (.ZN (n_0_0_87), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_441)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_245 (.ZN (n_0_250), .A (n_0_0_86));
AOI221_X1 i_0_0_244 (.ZN (n_0_0_86), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_442)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_243 (.ZN (n_0_249), .A (n_0_0_85));
AOI221_X1 i_0_0_242 (.ZN (n_0_0_85), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_443)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_241 (.ZN (n_0_248), .A (n_0_0_84));
AOI221_X1 i_0_0_240 (.ZN (n_0_0_84), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_444)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_239 (.ZN (n_0_247), .A (n_0_0_83));
AOI221_X1 i_0_0_238 (.ZN (n_0_0_83), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_445)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_237 (.ZN (n_0_246), .A (n_0_0_82));
AOI221_X1 i_0_0_236 (.ZN (n_0_0_82), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_446)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_235 (.ZN (n_0_245), .A (n_0_0_81));
AOI221_X1 i_0_0_234 (.ZN (n_0_0_81), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_447)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_233 (.ZN (n_0_244), .A (n_0_0_80));
AOI221_X1 i_0_0_232 (.ZN (n_0_0_80), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_448)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_231 (.ZN (n_0_243), .A (n_0_0_79));
AOI221_X1 i_0_0_230 (.ZN (n_0_0_79), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_449)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_229 (.ZN (n_0_242), .A (n_0_0_78));
AOI221_X1 i_0_0_228 (.ZN (n_0_0_78), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_450)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_227 (.ZN (n_0_241), .A (n_0_0_77));
AOI221_X1 i_0_0_226 (.ZN (n_0_0_77), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_451)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_225 (.ZN (n_0_240), .A (n_0_0_76));
AOI221_X1 i_0_0_224 (.ZN (n_0_0_76), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_452)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_223 (.ZN (n_0_239), .A (n_0_0_75));
AOI221_X1 i_0_0_222 (.ZN (n_0_0_75), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_453)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_221 (.ZN (n_0_238), .A (n_0_0_74));
AOI221_X1 i_0_0_220 (.ZN (n_0_0_74), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_454)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_219 (.ZN (n_0_237), .A (n_0_0_73));
AOI221_X1 i_0_0_218 (.ZN (n_0_0_73), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_455)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_217 (.ZN (n_0_236), .A (n_0_0_72));
AOI221_X1 i_0_0_216 (.ZN (n_0_0_72), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_456)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_215 (.ZN (n_0_235), .A (n_0_0_71));
AOI221_X1 i_0_0_214 (.ZN (n_0_0_71), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_457)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_213 (.ZN (n_0_234), .A (n_0_0_70));
AOI221_X1 i_0_0_212 (.ZN (n_0_0_70), .A (n_0_0_67), .B1 (hfn_ipo_n21), .B2 (n_0_458)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_211 (.ZN (n_0_233), .A (n_0_0_69));
AOI221_X1 i_0_0_210 (.ZN (n_0_0_69), .A (n_0_0_67), .B1 (hfn_ipo_n22), .B2 (n_0_459)
    , .C1 (hfn_ipo_n19), .C2 (n_0_71));
INV_X1 i_0_0_209 (.ZN (n_0_232), .A (n_0_0_68));
AOI221_X1 i_0_0_208 (.ZN (n_0_0_68), .A (n_0_0_67), .B1 (hfn_ipo_n22), .B2 (n_0_460)
    , .C1 (hfn_ipo_n20), .C2 (n_0_70));
AND2_X2 i_0_0_207 (.ZN (n_0_0_67), .A1 (n_0_0_35), .A2 (n_0_335));
INV_X1 i_0_0_206 (.ZN (n_0_231), .A (n_0_0_66));
AOI222_X1 i_0_0_205 (.ZN (n_0_0_66), .A1 (n_0_0_35), .A2 (n_0_334), .B1 (hfn_ipo_n22)
    , .B2 (n_0_461), .C1 (hfn_ipo_n20), .C2 (n_0_69));
INV_X1 i_0_0_204 (.ZN (n_0_230), .A (n_0_0_65));
AOI222_X1 i_0_0_203 (.ZN (n_0_0_65), .A1 (n_0_0_35), .A2 (n_0_333), .B1 (hfn_ipo_n22)
    , .B2 (n_0_462), .C1 (hfn_ipo_n20), .C2 (n_0_68));
INV_X1 i_0_0_202 (.ZN (n_0_229), .A (n_0_0_64));
AOI222_X1 i_0_0_201 (.ZN (n_0_0_64), .A1 (n_0_0_35), .A2 (n_0_332), .B1 (hfn_ipo_n22)
    , .B2 (n_0_463), .C1 (hfn_ipo_n20), .C2 (n_0_67));
INV_X1 i_0_0_200 (.ZN (n_0_228), .A (n_0_0_63));
AOI222_X1 i_0_0_199 (.ZN (n_0_0_63), .A1 (n_0_0_35), .A2 (n_0_331), .B1 (hfn_ipo_n22)
    , .B2 (n_0_464), .C1 (hfn_ipo_n20), .C2 (n_0_66));
INV_X1 i_0_0_198 (.ZN (n_0_227), .A (n_0_0_62));
AOI222_X1 i_0_0_197 (.ZN (n_0_0_62), .A1 (n_0_0_35), .A2 (n_0_330), .B1 (hfn_ipo_n22)
    , .B2 (n_0_465), .C1 (hfn_ipo_n20), .C2 (n_0_65));
INV_X1 i_0_0_196 (.ZN (n_0_226), .A (n_0_0_61));
AOI222_X1 i_0_0_195 (.ZN (n_0_0_61), .A1 (n_0_0_35), .A2 (n_0_329), .B1 (hfn_ipo_n22)
    , .B2 (n_0_466), .C1 (hfn_ipo_n20), .C2 (n_0_64));
INV_X1 i_0_0_194 (.ZN (n_0_225), .A (n_0_0_60));
AOI222_X1 i_0_0_193 (.ZN (n_0_0_60), .A1 (n_0_0_35), .A2 (n_0_328), .B1 (hfn_ipo_n22)
    , .B2 (n_0_467), .C1 (hfn_ipo_n20), .C2 (n_0_63));
INV_X1 i_0_0_192 (.ZN (n_0_224), .A (n_0_0_59));
AOI222_X1 i_0_0_191 (.ZN (n_0_0_59), .A1 (n_0_0_35), .A2 (n_0_327), .B1 (hfn_ipo_n22)
    , .B2 (n_0_468), .C1 (hfn_ipo_n20), .C2 (n_0_62));
INV_X1 i_0_0_190 (.ZN (n_0_223), .A (n_0_0_58));
AOI222_X1 i_0_0_189 (.ZN (n_0_0_58), .A1 (n_0_0_35), .A2 (n_0_326), .B1 (hfn_ipo_n22)
    , .B2 (n_0_469), .C1 (hfn_ipo_n20), .C2 (n_0_61));
INV_X1 i_0_0_188 (.ZN (n_0_222), .A (n_0_0_57));
AOI222_X1 i_0_0_187 (.ZN (n_0_0_57), .A1 (n_0_0_35), .A2 (n_0_325), .B1 (hfn_ipo_n22)
    , .B2 (n_0_470), .C1 (hfn_ipo_n20), .C2 (n_0_60));
INV_X1 i_0_0_186 (.ZN (n_0_221), .A (n_0_0_56));
AOI222_X1 i_0_0_185 (.ZN (n_0_0_56), .A1 (n_0_0_35), .A2 (n_0_324), .B1 (hfn_ipo_n22)
    , .B2 (n_0_471), .C1 (hfn_ipo_n20), .C2 (n_0_59));
INV_X1 i_0_0_184 (.ZN (n_0_220), .A (n_0_0_55));
AOI222_X1 i_0_0_183 (.ZN (n_0_0_55), .A1 (n_0_0_35), .A2 (n_0_323), .B1 (hfn_ipo_n22)
    , .B2 (n_0_472), .C1 (hfn_ipo_n20), .C2 (n_0_58));
INV_X1 i_0_0_182 (.ZN (n_0_219), .A (n_0_0_54));
AOI222_X1 i_0_0_181 (.ZN (n_0_0_54), .A1 (n_0_0_35), .A2 (n_0_322), .B1 (hfn_ipo_n22)
    , .B2 (n_0_473), .C1 (hfn_ipo_n20), .C2 (n_0_57));
INV_X1 i_0_0_180 (.ZN (n_0_218), .A (n_0_0_53));
AOI222_X1 i_0_0_179 (.ZN (n_0_0_53), .A1 (n_0_0_35), .A2 (n_0_321), .B1 (hfn_ipo_n22)
    , .B2 (n_0_474), .C1 (hfn_ipo_n20), .C2 (n_0_56));
INV_X1 i_0_0_178 (.ZN (n_0_217), .A (n_0_0_52));
AOI222_X1 i_0_0_177 (.ZN (n_0_0_52), .A1 (n_0_0_35), .A2 (n_0_320), .B1 (hfn_ipo_n22)
    , .B2 (n_0_475), .C1 (hfn_ipo_n20), .C2 (n_0_55));
INV_X1 i_0_0_176 (.ZN (n_0_216), .A (n_0_0_51));
AOI222_X1 i_0_0_175 (.ZN (n_0_0_51), .A1 (n_0_0_35), .A2 (n_0_319), .B1 (hfn_ipo_n22)
    , .B2 (n_0_476), .C1 (hfn_ipo_n20), .C2 (n_0_54));
INV_X1 i_0_0_174 (.ZN (n_0_215), .A (n_0_0_50));
AOI222_X1 i_0_0_173 (.ZN (n_0_0_50), .A1 (n_0_0_35), .A2 (n_0_318), .B1 (hfn_ipo_n22)
    , .B2 (n_0_477), .C1 (hfn_ipo_n20), .C2 (n_0_53));
INV_X1 i_0_0_172 (.ZN (n_0_214), .A (n_0_0_49));
AOI222_X1 i_0_0_171 (.ZN (n_0_0_49), .A1 (n_0_0_35), .A2 (n_0_317), .B1 (hfn_ipo_n22)
    , .B2 (n_0_478), .C1 (hfn_ipo_n20), .C2 (n_0_52));
INV_X1 i_0_0_170 (.ZN (n_0_213), .A (n_0_0_48));
AOI222_X1 i_0_0_169 (.ZN (n_0_0_48), .A1 (n_0_0_35), .A2 (n_0_316), .B1 (hfn_ipo_n22)
    , .B2 (n_0_479), .C1 (hfn_ipo_n20), .C2 (n_0_51));
INV_X1 i_0_0_168 (.ZN (n_0_212), .A (n_0_0_47));
AOI222_X1 i_0_0_167 (.ZN (n_0_0_47), .A1 (n_0_0_35), .A2 (n_0_315), .B1 (hfn_ipo_n22)
    , .B2 (n_0_480), .C1 (hfn_ipo_n20), .C2 (n_0_50));
INV_X1 i_0_0_166 (.ZN (n_0_211), .A (n_0_0_46));
AOI222_X1 i_0_0_165 (.ZN (n_0_0_46), .A1 (n_0_0_35), .A2 (n_0_314), .B1 (hfn_ipo_n22)
    , .B2 (n_0_481), .C1 (hfn_ipo_n20), .C2 (n_0_49));
INV_X1 i_0_0_164 (.ZN (n_0_210), .A (n_0_0_45));
AOI222_X1 i_0_0_163 (.ZN (n_0_0_45), .A1 (n_0_0_35), .A2 (n_0_313), .B1 (hfn_ipo_n22)
    , .B2 (n_0_482), .C1 (hfn_ipo_n20), .C2 (n_0_48));
INV_X1 i_0_0_162 (.ZN (n_0_209), .A (n_0_0_44));
AOI222_X1 i_0_0_161 (.ZN (n_0_0_44), .A1 (n_0_0_35), .A2 (n_0_312), .B1 (hfn_ipo_n22)
    , .B2 (n_0_483), .C1 (hfn_ipo_n19), .C2 (n_0_47));
INV_X1 i_0_0_160 (.ZN (n_0_208), .A (n_0_0_43));
AOI222_X1 i_0_0_159 (.ZN (n_0_0_43), .A1 (n_0_0_35), .A2 (n_0_311), .B1 (hfn_ipo_n21)
    , .B2 (n_0_484), .C1 (hfn_ipo_n19), .C2 (n_0_46));
INV_X1 i_0_0_158 (.ZN (n_0_207), .A (n_0_0_42));
AOI222_X1 i_0_0_157 (.ZN (n_0_0_42), .A1 (n_0_0_35), .A2 (n_0_310), .B1 (hfn_ipo_n21)
    , .B2 (n_0_485), .C1 (hfn_ipo_n19), .C2 (n_0_45));
INV_X1 i_0_0_156 (.ZN (n_0_206), .A (n_0_0_41));
AOI222_X1 i_0_0_155 (.ZN (n_0_0_41), .A1 (n_0_0_35), .A2 (n_0_309), .B1 (hfn_ipo_n21)
    , .B2 (n_0_486), .C1 (hfn_ipo_n19), .C2 (n_0_44));
INV_X1 i_0_0_154 (.ZN (n_0_205), .A (n_0_0_40));
AOI222_X1 i_0_0_153 (.ZN (n_0_0_40), .A1 (n_0_0_35), .A2 (n_0_308), .B1 (hfn_ipo_n22)
    , .B2 (n_0_487), .C1 (hfn_ipo_n20), .C2 (n_0_43));
INV_X1 i_0_0_152 (.ZN (n_0_204), .A (n_0_0_39));
AOI222_X1 i_0_0_151 (.ZN (n_0_0_39), .A1 (n_0_0_35), .A2 (n_0_307), .B1 (hfn_ipo_n22)
    , .B2 (n_0_488), .C1 (hfn_ipo_n20), .C2 (n_0_42));
INV_X1 i_0_0_150 (.ZN (n_0_203), .A (n_0_0_38));
AOI222_X1 i_0_0_149 (.ZN (n_0_0_38), .A1 (n_0_0_35), .A2 (n_0_306), .B1 (hfn_ipo_n22)
    , .B2 (n_0_489), .C1 (hfn_ipo_n20), .C2 (n_0_41));
INV_X1 i_0_0_148 (.ZN (n_0_202), .A (n_0_0_37));
AOI222_X1 i_0_0_147 (.ZN (n_0_0_37), .A1 (n_0_0_35), .A2 (n_0_305), .B1 (hfn_ipo_n22)
    , .B2 (n_0_490), .C1 (hfn_ipo_n20), .C2 (n_0_40));
INV_X1 i_0_0_146 (.ZN (n_0_201), .A (n_0_0_101));
NOR2_X1 i_0_0_145 (.ZN (n_0_0_36), .A1 (hfn_ipo_n20), .A2 (drc_ipo_n89));
NOR2_X4 i_0_0_144 (.ZN (n_0_0_35), .A1 (hfn_ipo_n20), .A2 (n_0_0_103));
AND2_X1 i_0_0_143 (.ZN (n_0_0_34), .A1 (n_0_0_110), .A2 (drc_ipo_n89));
OR2_X1 i_0_0_142 (.ZN (n_0_265), .A1 (drc_ipo_n89), .A2 (n_0_0_102));
AND2_X1 i_0_0_141 (.ZN (n_0_271), .A1 (n_0_0_103), .A2 (n_0_0_109));
AND2_X1 i_0_0_140 (.ZN (n_0_270), .A1 (n_0_0_103), .A2 (n_0_0_108));
AND2_X1 i_0_0_139 (.ZN (n_0_269), .A1 (n_0_0_103), .A2 (n_0_0_107));
AND2_X1 i_0_0_138 (.ZN (n_0_268), .A1 (n_0_0_103), .A2 (n_0_0_106));
AND2_X1 i_0_0_137 (.ZN (n_0_267), .A1 (n_0_0_103), .A2 (n_0_0_105));
AND2_X1 i_0_0_136 (.ZN (n_0_266), .A1 (n_0_0_103), .A2 (n_0_0_104));
NAND2_X1 i_0_0_135 (.ZN (n_0_272), .A1 (n_0_0_112), .A2 (n_0_0_103));
NAND2_X1 i_0_0_134 (.ZN (n_0_0_112), .A1 (n_0_0_111), .A2 (n_0_0_102));
MUX2_X1 i_0_0_133 (.Z (n_0_0_111), .A (n_0_0_18), .B (n_0_0_33), .S (\ctr[4] ));
MUX2_X1 i_0_0_132 (.Z (n_0_0_33), .A (n_0_0_25), .B (n_0_0_32), .S (\ctr[3] ));
MUX2_X1 i_0_0_131 (.Z (n_0_0_32), .A (n_0_0_28), .B (n_0_0_31), .S (\ctr[2] ));
MUX2_X1 i_0_0_130 (.Z (n_0_0_31), .A (n_0_0_29), .B (n_0_0_30), .S (\ctr[1] ));
MUX2_X1 i_0_0_129 (.Z (n_0_0_30), .A (\multiplier[30] ), .B (\multiplier[31] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_128 (.Z (n_0_0_29), .A (\multiplier[28] ), .B (\multiplier[29] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_127 (.Z (n_0_0_28), .A (n_0_0_26), .B (n_0_0_27), .S (\ctr[1] ));
MUX2_X1 i_0_0_126 (.Z (n_0_0_27), .A (\multiplier[26] ), .B (\multiplier[27] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_125 (.Z (n_0_0_26), .A (\multiplier[24] ), .B (\multiplier[25] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_124 (.Z (n_0_0_25), .A (n_0_0_21), .B (n_0_0_24), .S (\ctr[2] ));
MUX2_X1 i_0_0_123 (.Z (n_0_0_24), .A (n_0_0_22), .B (n_0_0_23), .S (\ctr[1] ));
MUX2_X1 i_0_0_122 (.Z (n_0_0_23), .A (\multiplier[22] ), .B (\multiplier[23] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_121 (.Z (n_0_0_22), .A (\multiplier[20] ), .B (\multiplier[21] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_120 (.Z (n_0_0_21), .A (n_0_0_19), .B (n_0_0_20), .S (\ctr[1] ));
MUX2_X1 i_0_0_119 (.Z (n_0_0_20), .A (\multiplier[18] ), .B (\multiplier[19] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_118 (.Z (n_0_0_19), .A (\multiplier[16] ), .B (\multiplier[17] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_117 (.Z (n_0_0_18), .A (n_0_0_10), .B (n_0_0_17), .S (\ctr[3] ));
MUX2_X1 i_0_0_116 (.Z (n_0_0_17), .A (n_0_0_13), .B (n_0_0_16), .S (\ctr[2] ));
MUX2_X1 i_0_0_115 (.Z (n_0_0_16), .A (n_0_0_14), .B (n_0_0_15), .S (\ctr[1] ));
MUX2_X1 i_0_0_114 (.Z (n_0_0_15), .A (\multiplier[14] ), .B (\multiplier[15] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_113 (.Z (n_0_0_14), .A (\multiplier[12] ), .B (\multiplier[13] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_112 (.Z (n_0_0_13), .A (n_0_0_11), .B (n_0_0_12), .S (\ctr[1] ));
MUX2_X1 i_0_0_111 (.Z (n_0_0_12), .A (\multiplier[10] ), .B (\multiplier[11] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_110 (.Z (n_0_0_11), .A (\multiplier[8] ), .B (\multiplier[9] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_109 (.Z (n_0_0_10), .A (n_0_0_6), .B (n_0_0_9), .S (\ctr[2] ));
MUX2_X1 i_0_0_108 (.Z (n_0_0_9), .A (n_0_0_7), .B (n_0_0_8), .S (\ctr[1] ));
MUX2_X1 i_0_0_107 (.Z (n_0_0_8), .A (\multiplier[6] ), .B (\multiplier[7] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_106 (.Z (n_0_0_7), .A (\multiplier[4] ), .B (\multiplier[5] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_105 (.Z (n_0_0_6), .A (n_0_0_4), .B (n_0_0_5), .S (\ctr[1] ));
MUX2_X1 i_0_0_104 (.Z (n_0_0_5), .A (\multiplier[2] ), .B (\multiplier[3] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_103 (.Z (n_0_0_4), .A (\multiplier[0] ), .B (\multiplier[1] ), .S (\ctr[0] ));
MUX2_X1 i_0_0_102 (.Z (n_0_303), .A (n_0_39), .B (n_0_367), .S (n_0_0_113));
MUX2_X1 i_0_0_101 (.Z (n_0_302), .A (n_0_38), .B (n_0_366), .S (n_0_0_113));
MUX2_X1 i_0_0_100 (.Z (n_0_301), .A (n_0_37), .B (n_0_365), .S (n_0_0_113));
MUX2_X1 i_0_0_99 (.Z (n_0_300), .A (n_0_36), .B (n_0_364), .S (n_0_0_113));
MUX2_X1 i_0_0_98 (.Z (n_0_299), .A (n_0_35), .B (n_0_363), .S (n_0_0_113));
MUX2_X1 i_0_0_97 (.Z (n_0_298), .A (n_0_34), .B (n_0_362), .S (n_0_0_113));
MUX2_X1 i_0_0_96 (.Z (n_0_297), .A (n_0_33), .B (n_0_361), .S (n_0_0_113));
MUX2_X1 i_0_0_95 (.Z (n_0_296), .A (n_0_32), .B (n_0_360), .S (n_0_0_113));
MUX2_X1 i_0_0_94 (.Z (n_0_295), .A (n_0_31), .B (n_0_359), .S (n_0_0_113));
MUX2_X1 i_0_0_93 (.Z (n_0_294), .A (n_0_30), .B (n_0_358), .S (n_0_0_113));
MUX2_X1 i_0_0_92 (.Z (n_0_293), .A (n_0_29), .B (n_0_357), .S (n_0_0_113));
MUX2_X1 i_0_0_91 (.Z (n_0_292), .A (n_0_28), .B (n_0_356), .S (n_0_0_113));
MUX2_X1 i_0_0_90 (.Z (n_0_291), .A (n_0_27), .B (n_0_355), .S (n_0_0_113));
MUX2_X1 i_0_0_89 (.Z (n_0_290), .A (n_0_26), .B (n_0_354), .S (n_0_0_113));
MUX2_X1 i_0_0_88 (.Z (n_0_289), .A (n_0_25), .B (n_0_353), .S (n_0_0_113));
MUX2_X1 i_0_0_87 (.Z (n_0_288), .A (n_0_24), .B (n_0_352), .S (n_0_0_113));
MUX2_X1 i_0_0_86 (.Z (n_0_287), .A (n_0_23), .B (n_0_351), .S (n_0_0_113));
MUX2_X1 i_0_0_85 (.Z (n_0_286), .A (n_0_22), .B (n_0_350), .S (n_0_0_113));
MUX2_X1 i_0_0_84 (.Z (n_0_285), .A (n_0_21), .B (n_0_349), .S (n_0_0_113));
MUX2_X1 i_0_0_83 (.Z (n_0_284), .A (n_0_20), .B (n_0_348), .S (n_0_0_113));
MUX2_X1 i_0_0_82 (.Z (n_0_283), .A (n_0_19), .B (n_0_347), .S (n_0_0_113));
MUX2_X1 i_0_0_81 (.Z (n_0_282), .A (n_0_18), .B (n_0_346), .S (n_0_0_113));
MUX2_X1 i_0_0_80 (.Z (n_0_281), .A (n_0_17), .B (n_0_345), .S (n_0_0_113));
MUX2_X1 i_0_0_79 (.Z (n_0_280), .A (n_0_16), .B (n_0_344), .S (n_0_0_113));
MUX2_X1 i_0_0_78 (.Z (n_0_279), .A (n_0_15), .B (n_0_343), .S (n_0_0_113));
MUX2_X1 i_0_0_77 (.Z (n_0_278), .A (n_0_14), .B (n_0_342), .S (n_0_0_113));
MUX2_X1 i_0_0_76 (.Z (n_0_277), .A (n_0_13), .B (n_0_341), .S (n_0_0_113));
MUX2_X1 i_0_0_75 (.Z (n_0_276), .A (n_0_12), .B (n_0_340), .S (n_0_0_113));
MUX2_X1 i_0_0_74 (.Z (n_0_275), .A (n_0_11), .B (n_0_339), .S (n_0_0_113));
MUX2_X1 i_0_0_73 (.Z (n_0_274), .A (n_0_10), .B (n_0_338), .S (n_0_0_113));
MUX2_X1 i_0_0_72 (.Z (n_0_273), .A (n_0_9), .B (n_0_337), .S (n_0_0_113));
AND2_X1 i_0_0_71 (.ZN (n_0_0_110), .A1 (n_0_367), .A2 (n_0_335));
OR2_X1 i_0_0_70 (.ZN (n_0_335), .A1 (drc_ipo_n56), .A2 (hfn_ipo_n18));
MUX2_X1 i_0_0_69 (.Z (n_0_334), .A (drc_ipo_n55), .B (drc_ipo_n87), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_68 (.Z (n_0_333), .A (drc_ipo_n54), .B (drc_ipo_n86), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_67 (.Z (n_0_332), .A (drc_ipo_n53), .B (drc_ipo_n85), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_66 (.Z (n_0_331), .A (drc_ipo_n52), .B (drc_ipo_n84), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_65 (.Z (n_0_330), .A (drc_ipo_n51), .B (drc_ipo_n83), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_64 (.Z (n_0_329), .A (drc_ipo_n50), .B (drc_ipo_n82), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_63 (.Z (n_0_328), .A (drc_ipo_n49), .B (drc_ipo_n81), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_62 (.Z (n_0_327), .A (drc_ipo_n48), .B (drc_ipo_n80), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_61 (.Z (n_0_326), .A (drc_ipo_n47), .B (drc_ipo_n79), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_60 (.Z (n_0_325), .A (drc_ipo_n46), .B (drc_ipo_n78), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_59 (.Z (n_0_324), .A (drc_ipo_n45), .B (drc_ipo_n77), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_58 (.Z (n_0_323), .A (drc_ipo_n44), .B (drc_ipo_n76), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_57 (.Z (n_0_322), .A (drc_ipo_n43), .B (drc_ipo_n75), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_56 (.Z (n_0_321), .A (drc_ipo_n42), .B (drc_ipo_n74), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_55 (.Z (n_0_320), .A (drc_ipo_n41), .B (drc_ipo_n73), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_54 (.Z (n_0_319), .A (drc_ipo_n40), .B (drc_ipo_n72), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_53 (.Z (n_0_318), .A (drc_ipo_n39), .B (drc_ipo_n71), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_52 (.Z (n_0_317), .A (drc_ipo_n38), .B (drc_ipo_n70), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_51 (.Z (n_0_316), .A (drc_ipo_n37), .B (drc_ipo_n69), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_50 (.Z (n_0_315), .A (drc_ipo_n36), .B (drc_ipo_n68), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_49 (.Z (n_0_314), .A (drc_ipo_n35), .B (drc_ipo_n67), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_48 (.Z (n_0_313), .A (drc_ipo_n34), .B (drc_ipo_n66), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_47 (.Z (n_0_312), .A (drc_ipo_n33), .B (drc_ipo_n65), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_46 (.Z (n_0_311), .A (drc_ipo_n32), .B (drc_ipo_n64), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_45 (.Z (n_0_310), .A (drc_ipo_n31), .B (drc_ipo_n63), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_44 (.Z (n_0_309), .A (drc_ipo_n30), .B (drc_ipo_n62), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_43 (.Z (n_0_308), .A (drc_ipo_n29), .B (drc_ipo_n61), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_42 (.Z (n_0_307), .A (drc_ipo_n28), .B (drc_ipo_n60), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_41 (.Z (n_0_306), .A (drc_ipo_n27), .B (drc_ipo_n59), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_40 (.Z (n_0_305), .A (drc_ipo_n26), .B (drc_ipo_n58), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_39 (.Z (n_0_304), .A (drc_ipo_n25), .B (drc_ipo_n57), .S (hfn_ipo_n17));
AND2_X1 i_0_0_38 (.ZN (n_0_367), .A1 (drc_ipo_n56), .A2 (hfn_ipo_n18));
MUX2_X1 i_0_0_37 (.Z (n_0_366), .A (drc_ipo_n87), .B (drc_ipo_n55), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_36 (.Z (n_0_365), .A (drc_ipo_n86), .B (drc_ipo_n54), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_35 (.Z (n_0_364), .A (drc_ipo_n85), .B (drc_ipo_n53), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_34 (.Z (n_0_363), .A (drc_ipo_n84), .B (drc_ipo_n52), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_33 (.Z (n_0_362), .A (drc_ipo_n83), .B (drc_ipo_n51), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_32 (.Z (n_0_361), .A (drc_ipo_n82), .B (drc_ipo_n50), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_31 (.Z (n_0_360), .A (drc_ipo_n81), .B (drc_ipo_n49), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_30 (.Z (n_0_359), .A (drc_ipo_n80), .B (drc_ipo_n48), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_29 (.Z (n_0_358), .A (drc_ipo_n79), .B (drc_ipo_n47), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_28 (.Z (n_0_357), .A (drc_ipo_n78), .B (drc_ipo_n46), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_27 (.Z (n_0_356), .A (drc_ipo_n77), .B (drc_ipo_n45), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_26 (.Z (n_0_355), .A (drc_ipo_n76), .B (drc_ipo_n44), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_25 (.Z (n_0_354), .A (drc_ipo_n75), .B (drc_ipo_n43), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_24 (.Z (n_0_353), .A (drc_ipo_n74), .B (drc_ipo_n42), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_23 (.Z (n_0_352), .A (drc_ipo_n73), .B (drc_ipo_n41), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_22 (.Z (n_0_351), .A (drc_ipo_n72), .B (drc_ipo_n40), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_21 (.Z (n_0_350), .A (drc_ipo_n71), .B (drc_ipo_n39), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_20 (.Z (n_0_349), .A (drc_ipo_n70), .B (drc_ipo_n38), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_19 (.Z (n_0_348), .A (drc_ipo_n69), .B (drc_ipo_n37), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_18 (.Z (n_0_347), .A (drc_ipo_n68), .B (drc_ipo_n36), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_17 (.Z (n_0_346), .A (drc_ipo_n67), .B (drc_ipo_n35), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_16 (.Z (n_0_345), .A (drc_ipo_n66), .B (drc_ipo_n34), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_15 (.Z (n_0_344), .A (drc_ipo_n65), .B (drc_ipo_n33), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_14 (.Z (n_0_343), .A (drc_ipo_n64), .B (drc_ipo_n32), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_13 (.Z (n_0_342), .A (drc_ipo_n63), .B (drc_ipo_n31), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_12 (.Z (n_0_341), .A (drc_ipo_n62), .B (drc_ipo_n30), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_11 (.Z (n_0_340), .A (drc_ipo_n61), .B (drc_ipo_n29), .S (hfn_ipo_n18));
MUX2_X1 i_0_0_10 (.Z (n_0_339), .A (drc_ipo_n60), .B (drc_ipo_n28), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_9 (.Z (n_0_338), .A (drc_ipo_n59), .B (drc_ipo_n27), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_8 (.Z (n_0_337), .A (drc_ipo_n58), .B (drc_ipo_n26), .S (hfn_ipo_n17));
MUX2_X1 i_0_0_7 (.Z (n_0_336), .A (drc_ipo_n57), .B (drc_ipo_n25), .S (hfn_ipo_n17));
NOR4_X1 i_0_0_6 (.ZN (n_0_368), .A1 (n_0_0_3), .A2 (\ctr[0] ), .A3 (\ctr[1] ), .A4 (\ctr[2] ));
OR4_X1 i_0_0_5 (.ZN (n_0_0_3), .A1 (n_0_0_102), .A2 (\ctr[3] ), .A3 (\ctr[4] ), .A4 (drc_ipo_n89));
HA_X1 i_0_0_4 (.CO (n_0_0_109), .S (n_0_0_108), .A (\ctr[4] ), .B (n_0_0_2));
HA_X1 i_0_0_3 (.CO (n_0_0_2), .S (n_0_0_107), .A (\ctr[3] ), .B (n_0_0_1));
HA_X1 i_0_0_2 (.CO (n_0_0_1), .S (n_0_0_106), .A (\ctr[2] ), .B (n_0_0_0));
HA_X1 i_0_0_1 (.CO (n_0_0_0), .S (n_0_0_105), .A (\ctr[1] ), .B (\ctr[0] ));
INV_X1 i_0_0_0 (.ZN (n_0_0_104), .A (\ctr[0] ));
datapath__0_12 i_0_15 (.p_0 ({n_0_136, n_0_135, n_0_134, n_0_133, n_0_131, n_0_130, 
    n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, 
    n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
    n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, 
    n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, 
    n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, 
    n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, 
    n_0_72}), .accumulator ({n_0_372, n_0_373, n_0_374, n_0_375, n_0_376, n_0_377, 
    n_0_378, n_0_379, n_0_380, n_0_381, n_0_382, n_0_383, n_0_384, n_0_385, n_0_386, 
    n_0_387, n_0_388, n_0_389, n_0_390, n_0_391, n_0_392, n_0_393, n_0_394, n_0_395, 
    n_0_396, n_0_397, n_0_398, n_0_399, n_0_400, n_0_401, n_0_402, n_0_403, n_0_404, 
    n_0_405, n_0_406, n_0_407, n_0_408, n_0_409, n_0_410, n_0_411, n_0_412, n_0_413, 
    n_0_414, n_0_415, n_0_416, n_0_417, n_0_418, n_0_419, n_0_420, n_0_421, n_0_422, 
    n_0_423, n_0_424, n_0_425, n_0_426, n_0_427, n_0_1, n_0_2, n_0_3, n_0_4, n_0_5, 
    n_0_6, n_0_7, n_0_8}), .multiplicand ({n_0_369, n_0_428, n_0_429, n_0_430, n_0_431, 
    n_0_432, n_0_433, n_0_434, n_0_435, n_0_436, n_0_437, n_0_438, n_0_439, n_0_440, 
    n_0_441, n_0_442, n_0_443, n_0_444, n_0_445, n_0_446, n_0_447, n_0_448, n_0_449, 
    n_0_450, n_0_451, n_0_452, n_0_453, n_0_454, n_0_455, n_0_456, n_0_457, n_0_458, 
    n_0_459, n_0_460, n_0_461, n_0_462, n_0_463, n_0_464, n_0_465, n_0_466, n_0_467, 
    n_0_468, n_0_469, n_0_470, n_0_471, n_0_472, n_0_473, n_0_474, n_0_475, n_0_476, 
    n_0_477, n_0_478, n_0_479, n_0_480, n_0_481, n_0_482, n_0_483, n_0_484, n_0_485, 
    n_0_486, n_0_487, n_0_488, n_0_489, n_0_490}));
datapath__0_10 i_0_13 (.p_0 ({n_0_71, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
    uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, 
    uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, 
    n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, 
    n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, 
    n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, 
    n_0_40, uc_32}), .p_1 ({uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, 
    uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, 
    uc_52, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, 
    uc_63, uc_64, n_0_335, n_0_334, n_0_333, n_0_332, n_0_331, n_0_330, n_0_329, 
    n_0_328, n_0_327, n_0_326, n_0_325, n_0_324, n_0_323, n_0_322, n_0_321, n_0_320, 
    n_0_319, n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, n_0_311, 
    n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304}));
datapath i_0_3 (.p_0 ({n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, 
    n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, 
    n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, 
    n_0_11, n_0_10, n_0_9, uc_0}), .p_1 ({n_0_367, n_0_366, n_0_365, n_0_364, n_0_363, 
    n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, n_0_356, n_0_355, n_0_354, 
    n_0_353, n_0_352, n_0_351, n_0_350, n_0_349, n_0_348, n_0_347, n_0_346, n_0_345, 
    n_0_344, n_0_343, n_0_342, n_0_341, n_0_340, n_0_339, n_0_338, n_0_337, n_0_336}));
DFF_X1 \product_reg[0]  (.Q (product[0]), .CK (CTS_n_tid0_299), .D (n_0_8));
DFF_X1 \product_reg[1]  (.Q (product[1]), .CK (CTS_n_tid0_299), .D (n_0_7));
DFF_X1 \product_reg[2]  (.Q (product[2]), .CK (CTS_n_tid0_299), .D (n_0_6));
DFF_X1 \product_reg[3]  (.Q (product[3]), .CK (CTS_n_tid0_299), .D (n_0_5));
DFF_X1 \product_reg[4]  (.Q (product[4]), .CK (CTS_n_tid0_299), .D (n_0_4));
DFF_X1 \product_reg[5]  (.Q (product[5]), .CK (CTS_n_tid0_299), .D (n_0_3));
DFF_X1 \product_reg[6]  (.Q (product[6]), .CK (CTS_n_tid0_299), .D (n_0_2));
DFF_X1 \product_reg[7]  (.Q (product[7]), .CK (CTS_n_tid0_299), .D (n_0_1));
DFF_X1 \product_reg[8]  (.Q (product[8]), .CK (CTS_n_tid0_299), .D (n_0_427));
DFF_X1 \product_reg[9]  (.Q (product[9]), .CK (CTS_n_tid0_299), .D (n_0_426));
DFF_X1 \product_reg[10]  (.Q (product[10]), .CK (CTS_n_tid0_299), .D (n_0_425));
DFF_X1 \product_reg[11]  (.Q (product[11]), .CK (CTS_n_tid0_299), .D (n_0_424));
DFF_X1 \product_reg[12]  (.Q (product[12]), .CK (CTS_n_tid0_299), .D (n_0_423));
DFF_X1 \product_reg[13]  (.Q (product[13]), .CK (CTS_n_tid0_299), .D (n_0_422));
DFF_X1 \product_reg[14]  (.Q (product[14]), .CK (CTS_n_tid0_299), .D (n_0_421));
DFF_X1 \product_reg[15]  (.Q (product[15]), .CK (CTS_n_tid0_299), .D (n_0_420));
DFF_X1 \product_reg[16]  (.Q (product[16]), .CK (CTS_n_tid0_299), .D (n_0_419));
DFF_X1 \product_reg[17]  (.Q (product[17]), .CK (CTS_n_tid0_299), .D (n_0_418));
DFF_X1 \product_reg[18]  (.Q (product[18]), .CK (CTS_n_tid0_299), .D (n_0_417));
DFF_X1 \product_reg[19]  (.Q (product[19]), .CK (CTS_n_tid0_299), .D (n_0_416));
DFF_X1 \product_reg[20]  (.Q (product[20]), .CK (CTS_n_tid0_299), .D (n_0_415));
DFF_X1 \product_reg[21]  (.Q (product[21]), .CK (CTS_n_tid0_299), .D (n_0_414));
DFF_X1 \product_reg[22]  (.Q (product[22]), .CK (CTS_n_tid0_299), .D (n_0_413));
DFF_X1 \product_reg[23]  (.Q (product[23]), .CK (CTS_n_tid0_299), .D (n_0_412));
DFF_X1 \product_reg[24]  (.Q (product[24]), .CK (CTS_n_tid0_299), .D (n_0_411));
DFF_X1 \product_reg[25]  (.Q (product[25]), .CK (CTS_n_tid0_299), .D (n_0_410));
DFF_X1 \product_reg[26]  (.Q (product[26]), .CK (CTS_n_tid0_299), .D (n_0_409));
DFF_X1 \product_reg[27]  (.Q (product[27]), .CK (CTS_n_tid0_299), .D (n_0_408));
DFF_X1 \product_reg[28]  (.Q (product[28]), .CK (CTS_n_tid0_299), .D (n_0_407));
DFF_X1 \product_reg[29]  (.Q (product[29]), .CK (CTS_n_tid0_299), .D (n_0_406));
DFF_X1 \product_reg[30]  (.Q (product[30]), .CK (CTS_n_tid0_299), .D (n_0_405));
DFF_X1 \product_reg[31]  (.Q (product[31]), .CK (CTS_n_tid0_299), .D (n_0_404));
DFF_X1 \product_reg[32]  (.Q (product[32]), .CK (CTS_n_tid0_299), .D (n_0_403));
DFF_X1 \product_reg[33]  (.Q (product[33]), .CK (CTS_n_tid0_299), .D (n_0_402));
DFF_X1 \product_reg[34]  (.Q (product[34]), .CK (CTS_n_tid0_299), .D (n_0_401));
DFF_X1 \product_reg[35]  (.Q (product[35]), .CK (CTS_n_tid0_299), .D (n_0_400));
DFF_X1 \product_reg[36]  (.Q (product[36]), .CK (CTS_n_tid0_299), .D (n_0_399));
DFF_X1 \product_reg[37]  (.Q (product[37]), .CK (CTS_n_tid0_299), .D (n_0_398));
DFF_X1 \product_reg[38]  (.Q (product[38]), .CK (CTS_n_tid0_299), .D (n_0_397));
DFF_X1 \product_reg[39]  (.Q (product[39]), .CK (CTS_n_tid0_299), .D (n_0_396));
DFF_X1 \product_reg[40]  (.Q (product[40]), .CK (CTS_n_tid0_299), .D (n_0_395));
DFF_X1 \product_reg[41]  (.Q (product[41]), .CK (CTS_n_tid0_299), .D (n_0_394));
DFF_X1 \product_reg[42]  (.Q (product[42]), .CK (CTS_n_tid0_299), .D (n_0_393));
DFF_X1 \product_reg[43]  (.Q (product[43]), .CK (CTS_n_tid0_299), .D (n_0_392));
DFF_X1 \product_reg[44]  (.Q (product[44]), .CK (CTS_n_tid0_299), .D (n_0_391));
DFF_X1 \product_reg[45]  (.Q (product[45]), .CK (CTS_n_tid0_299), .D (n_0_390));
DFF_X1 \product_reg[46]  (.Q (product[46]), .CK (CTS_n_tid0_299), .D (n_0_389));
DFF_X1 \product_reg[47]  (.Q (product[47]), .CK (CTS_n_tid0_299), .D (n_0_388));
DFF_X1 \product_reg[48]  (.Q (product[48]), .CK (CTS_n_tid0_299), .D (n_0_387));
DFF_X1 \product_reg[49]  (.Q (product[49]), .CK (CTS_n_tid0_299), .D (n_0_386));
DFF_X1 \product_reg[50]  (.Q (product[50]), .CK (CTS_n_tid0_299), .D (n_0_385));
DFF_X1 \product_reg[51]  (.Q (product[51]), .CK (CTS_n_tid0_299), .D (n_0_384));
DFF_X1 \product_reg[52]  (.Q (product[52]), .CK (CTS_n_tid0_299), .D (n_0_383));
DFF_X1 \product_reg[53]  (.Q (product[53]), .CK (CTS_n_tid0_299), .D (n_0_382));
DFF_X1 \product_reg[54]  (.Q (product[54]), .CK (CTS_n_tid0_299), .D (n_0_381));
DFF_X1 \product_reg[55]  (.Q (product[55]), .CK (CTS_n_tid0_299), .D (n_0_380));
DFF_X1 \product_reg[56]  (.Q (product[56]), .CK (CTS_n_tid0_299), .D (n_0_379));
DFF_X1 \product_reg[57]  (.Q (product[57]), .CK (CTS_n_tid0_299), .D (n_0_378));
DFF_X1 \product_reg[58]  (.Q (product[58]), .CK (CTS_n_tid0_299), .D (n_0_377));
DFF_X1 \product_reg[59]  (.Q (product[59]), .CK (CTS_n_tid0_299), .D (n_0_376));
DFF_X1 \product_reg[60]  (.Q (product[60]), .CK (CTS_n_tid0_299), .D (n_0_375));
DFF_X1 \product_reg[61]  (.Q (product[61]), .CK (CTS_n_tid0_299), .D (n_0_374));
DFF_X1 \product_reg[62]  (.Q (product[62]), .CK (CTS_n_tid0_299), .D (n_0_373));
DFF_X1 \product_reg[63]  (.Q (product[63]), .CK (CTS_n_tid0_299), .D (n_0_372));
CLKGATETST_X8 clk_gate_product_reg (.GCK (CTS_n_tid0_300), .CK (CTS_n_tid1_362), .E (n_0_368), .SE (1'b0 ));
BUF_X2 hfn_ipo_c19 (.Z (hfn_ipo_n19), .A (n_0_0_34));
BUF_X4 hfn_ipo_c20 (.Z (hfn_ipo_n20), .A (n_0_0_34));
CLKBUF_X2 hfn_ipo_c21 (.Z (hfn_ipo_n21), .A (n_0_0_36));
CLKBUF_X2 hfn_ipo_c22 (.Z (hfn_ipo_n22), .A (n_0_0_36));
BUF_X2 hfn_ipo_c24 (.Z (hfn_ipo_n24), .A (n_0_0_103));
CLKBUF_X2 hfn_ipo_c17 (.Z (hfn_ipo_n17), .A (drc_ipo_n88));
CLKBUF_X2 hfn_ipo_c18 (.Z (hfn_ipo_n18), .A (drc_ipo_n88));
CLKBUF_X1 drc_ipo_c25 (.Z (drc_ipo_n25), .A (y[0]));
CLKBUF_X1 drc_ipo_c26 (.Z (drc_ipo_n26), .A (y[1]));
CLKBUF_X1 drc_ipo_c27 (.Z (drc_ipo_n27), .A (y[2]));
CLKBUF_X1 drc_ipo_c28 (.Z (drc_ipo_n28), .A (y[3]));
CLKBUF_X1 drc_ipo_c29 (.Z (drc_ipo_n29), .A (y[4]));
CLKBUF_X1 drc_ipo_c30 (.Z (drc_ipo_n30), .A (y[5]));
CLKBUF_X1 drc_ipo_c31 (.Z (drc_ipo_n31), .A (y[6]));
CLKBUF_X1 drc_ipo_c32 (.Z (drc_ipo_n32), .A (y[7]));
CLKBUF_X1 drc_ipo_c33 (.Z (drc_ipo_n33), .A (y[8]));
CLKBUF_X1 drc_ipo_c34 (.Z (drc_ipo_n34), .A (y[9]));
CLKBUF_X1 drc_ipo_c35 (.Z (drc_ipo_n35), .A (y[10]));
CLKBUF_X1 drc_ipo_c36 (.Z (drc_ipo_n36), .A (y[11]));
CLKBUF_X1 drc_ipo_c37 (.Z (drc_ipo_n37), .A (y[12]));
CLKBUF_X1 drc_ipo_c38 (.Z (drc_ipo_n38), .A (y[13]));
CLKBUF_X1 drc_ipo_c39 (.Z (drc_ipo_n39), .A (y[14]));
CLKBUF_X1 drc_ipo_c40 (.Z (drc_ipo_n40), .A (y[15]));
CLKBUF_X1 drc_ipo_c41 (.Z (drc_ipo_n41), .A (y[16]));
CLKBUF_X1 drc_ipo_c42 (.Z (drc_ipo_n42), .A (y[17]));
CLKBUF_X1 drc_ipo_c43 (.Z (drc_ipo_n43), .A (y[18]));
CLKBUF_X1 drc_ipo_c44 (.Z (drc_ipo_n44), .A (y[19]));
CLKBUF_X1 drc_ipo_c45 (.Z (drc_ipo_n45), .A (y[20]));
CLKBUF_X1 drc_ipo_c46 (.Z (drc_ipo_n46), .A (y[21]));
CLKBUF_X1 drc_ipo_c47 (.Z (drc_ipo_n47), .A (y[22]));
CLKBUF_X1 drc_ipo_c48 (.Z (drc_ipo_n48), .A (y[23]));
CLKBUF_X1 drc_ipo_c49 (.Z (drc_ipo_n49), .A (y[24]));
CLKBUF_X1 drc_ipo_c50 (.Z (drc_ipo_n50), .A (y[25]));
CLKBUF_X1 drc_ipo_c51 (.Z (drc_ipo_n51), .A (y[26]));
CLKBUF_X1 drc_ipo_c52 (.Z (drc_ipo_n52), .A (y[27]));
CLKBUF_X1 drc_ipo_c53 (.Z (drc_ipo_n53), .A (y[28]));
CLKBUF_X1 drc_ipo_c54 (.Z (drc_ipo_n54), .A (y[29]));
CLKBUF_X1 drc_ipo_c55 (.Z (drc_ipo_n55), .A (y[30]));
CLKBUF_X1 drc_ipo_c56 (.Z (drc_ipo_n56), .A (y[31]));
CLKBUF_X1 drc_ipo_c57 (.Z (drc_ipo_n57), .A (x[0]));
CLKBUF_X1 drc_ipo_c58 (.Z (drc_ipo_n58), .A (x[1]));
CLKBUF_X1 drc_ipo_c59 (.Z (drc_ipo_n59), .A (x[2]));
CLKBUF_X1 drc_ipo_c60 (.Z (drc_ipo_n60), .A (x[3]));
CLKBUF_X1 drc_ipo_c61 (.Z (drc_ipo_n61), .A (x[4]));
CLKBUF_X1 drc_ipo_c62 (.Z (drc_ipo_n62), .A (x[5]));
CLKBUF_X1 drc_ipo_c63 (.Z (drc_ipo_n63), .A (x[6]));
CLKBUF_X1 drc_ipo_c64 (.Z (drc_ipo_n64), .A (x[7]));
CLKBUF_X1 drc_ipo_c65 (.Z (drc_ipo_n65), .A (x[8]));
CLKBUF_X1 drc_ipo_c66 (.Z (drc_ipo_n66), .A (x[9]));
CLKBUF_X1 drc_ipo_c67 (.Z (drc_ipo_n67), .A (x[10]));
CLKBUF_X1 drc_ipo_c68 (.Z (drc_ipo_n68), .A (x[11]));
CLKBUF_X1 drc_ipo_c69 (.Z (drc_ipo_n69), .A (x[12]));
CLKBUF_X1 drc_ipo_c70 (.Z (drc_ipo_n70), .A (x[13]));
CLKBUF_X1 drc_ipo_c71 (.Z (drc_ipo_n71), .A (x[14]));
CLKBUF_X1 drc_ipo_c72 (.Z (drc_ipo_n72), .A (x[15]));
CLKBUF_X1 drc_ipo_c73 (.Z (drc_ipo_n73), .A (x[16]));
CLKBUF_X1 drc_ipo_c74 (.Z (drc_ipo_n74), .A (x[17]));
CLKBUF_X1 drc_ipo_c75 (.Z (drc_ipo_n75), .A (x[18]));
CLKBUF_X1 drc_ipo_c76 (.Z (drc_ipo_n76), .A (x[19]));
CLKBUF_X1 drc_ipo_c77 (.Z (drc_ipo_n77), .A (x[20]));
CLKBUF_X1 drc_ipo_c78 (.Z (drc_ipo_n78), .A (x[21]));
CLKBUF_X1 drc_ipo_c79 (.Z (drc_ipo_n79), .A (x[22]));
CLKBUF_X1 drc_ipo_c80 (.Z (drc_ipo_n80), .A (x[23]));
CLKBUF_X1 drc_ipo_c81 (.Z (drc_ipo_n81), .A (x[24]));
CLKBUF_X1 drc_ipo_c82 (.Z (drc_ipo_n82), .A (x[25]));
CLKBUF_X1 drc_ipo_c83 (.Z (drc_ipo_n83), .A (x[26]));
CLKBUF_X1 drc_ipo_c84 (.Z (drc_ipo_n84), .A (x[27]));
CLKBUF_X1 drc_ipo_c85 (.Z (drc_ipo_n85), .A (x[28]));
CLKBUF_X1 drc_ipo_c86 (.Z (drc_ipo_n86), .A (x[29]));
CLKBUF_X1 drc_ipo_c87 (.Z (drc_ipo_n87), .A (x[30]));
CLKBUF_X1 drc_ipo_c88 (.Z (drc_ipo_n88), .A (x[31]));
CLKBUF_X1 drc_ipo_c89 (.Z (drc_ipo_n89), .A (rst));
CLKBUF_X3 CTS_L3_c_tid1_131 (.Z (CTS_n_tid1_126), .A (CTS_n_tid1_130));
CLKBUF_X2 CTS_L3_c_tid0_133 (.Z (CTS_n_tid0_128), .A (CTS_n_tid0_285));
CLKBUF_X2 CTS_L3_c_tid0_134 (.Z (CTS_n_tid0_129), .A (CTS_n_tid0_285));
CLKBUF_X3 CTS_L3_c_tid0_136 (.Z (CTS_n_tid0_132), .A (CTS_n_tid0_285));
CLKBUF_X3 CTS_L3_c_tid0_137 (.Z (CTS_n_tid0_133), .A (CTS_n_tid0_285));
CLKBUF_X3 CTS_L3_c_tid0_306 (.Z (CTS_n_tid0_299), .A (CTS_n_tid0_300));
CLKBUF_X2 CTS_L1_c_tid1_350 (.Z (CTS_n_tid1_362), .A (clk));

endmodule //sequential_multiplier


