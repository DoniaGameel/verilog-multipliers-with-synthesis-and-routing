/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Jan  4 11:38:34 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2946952376 */

module Reg__0_17(in, clk, out);
   input [31:0]in;
   input clk;
   output [31:0]out;

   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module Reg__0_18(in, clk, out);
   input [31:0]in;
   input clk;
   output [31:0]out;

   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module datapath(B, A, Out);
   input [23:0]B;
   input [23:0]A;
   output [47:0]Out;

   INV_X1 i_0 (.A(n_20), .ZN(Out[0]));
   AOI22_X1 i_1 (.A1(A[0]), .A2(B[1]), .B1(B[0]), .B2(A[1]), .ZN(n_3));
   NOR2_X1 i_2 (.A1(n_19), .A2(n_3), .ZN(Out[1]));
   NAND2_X1 i_3 (.A1(A[2]), .A2(B[3]), .ZN(n_30));
   OR3_X1 i_4 (.A1(n_30), .A2(n_1534), .A3(n_29), .ZN(n_32));
   OAI22_X1 i_5 (.A1(n_1534), .A2(n_424), .B1(n_29), .B2(n_33), .ZN(n_34));
   NAND2_X1 i_6 (.A1(n_32), .A2(n_34), .ZN(n_35));
   NAND2_X1 i_7 (.A1(A[0]), .A2(B[4]), .ZN(n_36));
   XNOR2_X1 i_8 (.A(n_35), .B(n_36), .ZN(n_37));
   NAND3_X1 i_9 (.A1(n_25), .A2(A[4]), .A3(n_107), .ZN(n_38));
   NAND2_X1 i_10 (.A1(B[1]), .A2(A[4]), .ZN(n_39));
   INV_X1 i_11 (.A(n_39), .ZN(n_40));
   OAI21_X1 i_12 (.A(n_107), .B1(n_25), .B2(n_40), .ZN(n_41));
   INV_X1 i_13 (.A(n_41), .ZN(n_42));
   AOI22_X1 i_14 (.A1(B[0]), .A2(A[4]), .B1(B[1]), .B2(A[3]), .ZN(n_43));
   OAI21_X1 i_15 (.A(n_38), .B1(n_42), .B2(n_43), .ZN(n_44));
   AOI21_X1 i_16 (.A(n_66), .B1(n_150), .B2(n_64), .ZN(n_45));
   NAND2_X1 i_17 (.A1(n_44), .A2(n_45), .ZN(n_46));
   OAI21_X1 i_18 (.A(n_46), .B1(n_44), .B2(n_45), .ZN(n_47));
   XOR2_X1 i_19 (.A(n_37), .B(n_47), .Z(n_48));
   OAI21_X1 i_20 (.A(n_143), .B1(n_141), .B2(n_149), .ZN(n_49));
   XNOR2_X1 i_21 (.A(n_48), .B(n_49), .ZN(Out[4]));
   OAI21_X1 i_22 (.A(n_32), .B1(n_35), .B2(n_36), .ZN(n_50));
   XNOR2_X1 i_23 (.A(n_50), .B(n_41), .ZN(n_51));
   NAND2_X1 i_24 (.A1(B[0]), .A2(A[5]), .ZN(n_52));
   XNOR2_X1 i_25 (.A(n_39), .B(n_52), .ZN(n_53));
   NAND2_X1 i_26 (.A1(B[2]), .A2(A[3]), .ZN(n_54));
   XOR2_X1 i_27 (.A(n_53), .B(n_54), .Z(n_55));
   XOR2_X1 i_28 (.A(n_51), .B(n_55), .Z(n_56));
   NAND2_X1 i_29 (.A1(A[1]), .A2(B[4]), .ZN(n_57));
   XNOR2_X1 i_30 (.A(n_30), .B(n_57), .ZN(n_58));
   NAND2_X1 i_31 (.A1(A[0]), .A2(B[5]), .ZN(n_59));
   XNOR2_X1 i_32 (.A(n_58), .B(n_59), .ZN(n_60));
   XOR2_X1 i_33 (.A(n_60), .B(n_46), .Z(n_61));
   XNOR2_X1 i_34 (.A(n_56), .B(n_61), .ZN(n_62));
   AOI22_X1 i_35 (.A1(n_48), .A2(n_49), .B1(n_47), .B2(n_37), .ZN(n_63));
   XNOR2_X1 i_36 (.A(n_62), .B(n_63), .ZN(Out[5]));
   NOR2_X1 i_37 (.A1(n_28), .A2(n_170), .ZN(n_65));
   OAI33_X1 i_38 (.A1(n_53), .A2(n_29), .A3(n_99), .B1(n_39), .B2(n_28), 
      .B3(n_423), .ZN(n_67));
   XOR2_X1 i_39 (.A(n_65), .B(n_67), .Z(n_68));
   OAI22_X1 i_40 (.A1(n_58), .A2(n_59), .B1(n_30), .B2(n_57), .ZN(n_69));
   XNOR2_X1 i_41 (.A(n_68), .B(n_69), .ZN(n_70));
   NAND2_X1 i_42 (.A1(A[2]), .A2(B[5]), .ZN(n_71));
   NOR2_X1 i_43 (.A1(n_57), .A2(n_71), .ZN(n_72));
   AOI22_X1 i_44 (.A1(A[2]), .A2(B[4]), .B1(A[1]), .B2(B[5]), .ZN(n_73));
   NOR2_X1 i_45 (.A1(n_72), .A2(n_73), .ZN(n_74));
   NAND2_X1 i_46 (.A1(A[0]), .A2(B[6]), .ZN(n_75));
   XNOR2_X1 i_47 (.A(n_74), .B(n_75), .ZN(n_76));
   NAND2_X1 i_48 (.A1(B[2]), .A2(A[5]), .ZN(n_77));
   NOR2_X1 i_49 (.A1(n_39), .A2(n_77), .ZN(n_78));
   AOI22_X1 i_50 (.A1(B[2]), .A2(A[4]), .B1(B[1]), .B2(A[5]), .ZN(n_79));
   NOR2_X1 i_51 (.A1(n_78), .A2(n_79), .ZN(n_80));
   NOR2_X1 i_52 (.A1(n_424), .A2(n_99), .ZN(n_81));
   XOR2_X1 i_53 (.A(n_80), .B(n_81), .Z(n_82));
   NAND2_X1 i_54 (.A1(n_76), .A2(n_82), .ZN(n_83));
   OAI21_X1 i_55 (.A(n_83), .B1(n_76), .B2(n_82), .ZN(n_84));
   XNOR2_X1 i_56 (.A(n_70), .B(n_84), .ZN(n_85));
   AOI22_X1 i_57 (.A1(n_51), .A2(n_55), .B1(n_50), .B2(n_42), .ZN(n_86));
   OAI21_X1 i_58 (.A(n_86), .B1(n_46), .B2(n_60), .ZN(n_87));
   OR3_X1 i_59 (.A1(n_86), .A2(n_46), .A3(n_60), .ZN(n_88));
   NAND2_X1 i_60 (.A1(n_87), .A2(n_88), .ZN(n_89));
   XOR2_X1 i_61 (.A(n_85), .B(n_89), .Z(n_90));
   OAI22_X1 i_62 (.A1(n_62), .A2(n_63), .B1(n_56), .B2(n_61), .ZN(n_91));
   XNOR2_X1 i_63 (.A(n_90), .B(n_91), .ZN(Out[6]));
   AOI22_X1 i_64 (.A1(n_68), .A2(n_69), .B1(n_67), .B2(n_65), .ZN(n_92));
   INV_X1 i_65 (.A(n_92), .ZN(n_93));
   INV_X1 i_66 (.A(n_75), .ZN(n_94));
   AOI21_X1 i_67 (.A(n_72), .B1(n_74), .B2(n_94), .ZN(n_95));
   INV_X1 i_68 (.A(n_95), .ZN(n_96));
   OAI22_X1 i_69 (.A1(n_93), .A2(n_95), .B1(n_92), .B2(n_96), .ZN(n_97));
   AOI21_X1 i_70 (.A(n_78), .B1(n_80), .B2(n_81), .ZN(n_98));
   NAND2_X1 i_71 (.A1(B[1]), .A2(A[6]), .ZN(n_100));
   XNOR2_X1 i_72 (.A(n_421), .B(n_100), .ZN(n_101));
   XOR2_X1 i_73 (.A(n_98), .B(n_101), .Z(n_102));
   XOR2_X1 i_74 (.A(n_97), .B(n_102), .Z(n_103));
   OAI21_X1 i_75 (.A(n_83), .B1(n_70), .B2(n_84), .ZN(n_104));
   NAND2_X1 i_76 (.A1(n_103), .A2(n_104), .ZN(n_105));
   OAI21_X1 i_77 (.A(n_105), .B1(n_103), .B2(n_104), .ZN(n_106));
   NOR2_X1 i_78 (.A1(n_75), .A2(n_386), .ZN(n_108));
   AOI22_X1 i_79 (.A1(A[1]), .A2(B[6]), .B1(A[0]), .B2(B[7]), .ZN(n_109));
   NOR2_X1 i_80 (.A1(n_108), .A2(n_109), .ZN(n_110));
   XNOR2_X1 i_81 (.A(n_110), .B(n_71), .ZN(n_111));
   NAND2_X1 i_82 (.A1(B[4]), .A2(A[3]), .ZN(n_112));
   OR3_X1 i_83 (.A1(n_77), .A2(n_424), .A3(n_422), .ZN(n_114));
   OAI21_X1 i_84 (.A(n_77), .B1(n_424), .B2(n_422), .ZN(n_115));
   NAND2_X1 i_85 (.A1(n_114), .A2(n_115), .ZN(n_116));
   XOR2_X1 i_86 (.A(n_112), .B(n_116), .Z(n_117));
   XOR2_X1 i_87 (.A(n_111), .B(n_117), .Z(n_118));
   XNOR2_X1 i_88 (.A(n_88), .B(n_118), .ZN(n_119));
   XNOR2_X1 i_89 (.A(n_106), .B(n_119), .ZN(n_120));
   AOI22_X1 i_90 (.A1(n_90), .A2(n_91), .B1(n_85), .B2(n_89), .ZN(n_121));
   XOR2_X1 i_91 (.A(n_120), .B(n_121), .Z(Out[7]));
   INV_X1 i_92 (.A(n_106), .ZN(n_122));
   AOI22_X1 i_93 (.A1(n_120), .A2(n_121), .B1(n_122), .B2(n_119), .ZN(n_123));
   AOI22_X1 i_94 (.A1(n_97), .A2(n_102), .B1(n_93), .B2(n_96), .ZN(n_124));
   OAI21_X1 i_95 (.A(n_114), .B1(n_116), .B2(n_112), .ZN(n_125));
   INV_X1 i_96 (.A(n_71), .ZN(n_126));
   AOI21_X1 i_97 (.A(n_108), .B1(n_110), .B2(n_126), .ZN(n_127));
   XNOR2_X1 i_98 (.A(n_125), .B(n_127), .ZN(n_128));
   OAI22_X1 i_99 (.A1(n_98), .A2(n_101), .B1(n_421), .B2(n_100), .ZN(n_129));
   XNOR2_X1 i_100 (.A(n_128), .B(n_129), .ZN(n_130));
   XOR2_X1 i_101 (.A(n_124), .B(n_130), .Z(n_131));
   XNOR2_X1 i_102 (.A(n_131), .B(n_105), .ZN(n_132));
   INV_X1 i_103 (.A(n_88), .ZN(n_133));
   AOI22_X1 i_104 (.A1(n_133), .A2(n_118), .B1(n_111), .B2(n_117), .ZN(n_134));
   NAND2_X1 i_105 (.A1(A[2]), .A2(B[6]), .ZN(n_135));
   XNOR2_X1 i_106 (.A(n_386), .B(n_135), .ZN(n_136));
   NAND2_X1 i_107 (.A1(A[0]), .A2(B[8]), .ZN(n_137));
   XOR2_X1 i_108 (.A(n_136), .B(n_137), .Z(n_138));
   XOR2_X1 i_109 (.A(n_417), .B(n_416), .Z(n_144));
   XNOR2_X1 i_110 (.A(n_138), .B(n_144), .ZN(n_145));
   XOR2_X1 i_111 (.A(n_393), .B(n_392), .Z(n_152));
   XOR2_X1 i_112 (.A(n_145), .B(n_152), .Z(n_153));
   NOR2_X1 i_113 (.A1(n_134), .A2(n_153), .ZN(n_154));
   AOI21_X1 i_114 (.A(n_154), .B1(n_134), .B2(n_153), .ZN(n_155));
   NAND2_X1 i_115 (.A1(n_132), .A2(n_155), .ZN(n_156));
   INV_X1 i_116 (.A(n_156), .ZN(n_157));
   NOR2_X1 i_117 (.A1(n_132), .A2(n_155), .ZN(n_158));
   NOR2_X1 i_118 (.A1(n_157), .A2(n_158), .ZN(n_159));
   XNOR2_X1 i_119 (.A(n_123), .B(n_159), .ZN(Out[8]));
   AOI21_X1 i_120 (.A(n_158), .B1(n_123), .B2(n_156), .ZN(n_160));
   AOI22_X1 i_121 (.A1(n_131), .A2(n_105), .B1(n_124), .B2(n_130), .ZN(n_161));
   NAND2_X1 i_122 (.A1(n_161), .A2(n_154), .ZN(n_162));
   OAI21_X1 i_123 (.A(n_162), .B1(n_161), .B2(n_154), .ZN(n_163));
   INV_X1 i_124 (.A(n_127), .ZN(n_164));
   AOI22_X1 i_125 (.A1(n_128), .A2(n_129), .B1(n_125), .B2(n_164), .ZN(n_165));
   XOR2_X1 i_126 (.A(n_381), .B(n_380), .Z(n_172));
   XOR2_X1 i_127 (.A(n_165), .B(n_172), .Z(n_173));
   XOR2_X1 i_128 (.A(n_397), .B(n_391), .Z(n_179));
   XOR2_X1 i_129 (.A(n_173), .B(n_179), .Z(n_180));
   NAND2_X1 i_130 (.A1(B[3]), .A2(A[6]), .ZN(n_183));
   XOR2_X1 i_131 (.A(n_454), .B(n_183), .Z(n_184));
   OAI22_X1 i_132 (.A1(n_136), .A2(n_137), .B1(n_386), .B2(n_135), .ZN(n_185));
   XOR2_X1 i_133 (.A(n_184), .B(n_185), .Z(n_186));
   XOR2_X1 i_134 (.A(n_388), .B(n_387), .Z(n_190));
   XNOR2_X1 i_135 (.A(n_186), .B(n_190), .ZN(n_191));
   OAI22_X1 i_136 (.A1(n_145), .A2(n_152), .B1(n_144), .B2(n_138), .ZN(n_192));
   NAND2_X1 i_137 (.A1(n_191), .A2(n_192), .ZN(n_193));
   OAI21_X1 i_138 (.A(n_193), .B1(n_191), .B2(n_192), .ZN(n_194));
   XNOR2_X1 i_139 (.A(n_180), .B(n_194), .ZN(n_195));
   NAND2_X1 i_140 (.A1(n_163), .A2(n_195), .ZN(n_196));
   OAI21_X1 i_141 (.A(n_196), .B1(n_163), .B2(n_195), .ZN(n_197));
   XNOR2_X1 i_142 (.A(n_160), .B(n_197), .ZN(Out[9]));
   NOR2_X1 i_143 (.A1(n_455), .A2(n_331), .ZN(n_199));
   AOI22_X1 i_144 (.A1(B[3]), .A2(A[7]), .B1(B[2]), .B2(A[8]), .ZN(n_200));
   NOR2_X1 i_145 (.A1(n_199), .A2(n_200), .ZN(n_201));
   NOR2_X1 i_146 (.A1(n_340), .A2(n_170), .ZN(n_202));
   XOR2_X1 i_147 (.A(n_201), .B(n_202), .Z(n_203));
   XOR2_X1 i_148 (.A(n_446), .B(n_445), .Z(n_210));
   XOR2_X1 i_149 (.A(n_203), .B(n_210), .Z(n_211));
   NAND2_X1 i_150 (.A1(B[5]), .A2(A[5]), .ZN(n_213));
   XNOR2_X1 i_151 (.A(n_370), .B(n_213), .ZN(n_214));
   NAND2_X1 i_152 (.A1(A[3]), .A2(B[7]), .ZN(n_215));
   XOR2_X1 i_153 (.A(n_214), .B(n_215), .Z(n_216));
   XNOR2_X1 i_154 (.A(n_211), .B(n_216), .ZN(n_217));
   INV_X1 i_155 (.A(n_165), .ZN(n_218));
   OAI22_X1 i_156 (.A1(n_173), .A2(n_179), .B1(n_218), .B2(n_172), .ZN(n_219));
   NAND2_X1 i_157 (.A1(n_217), .A2(n_219), .ZN(n_220));
   OAI21_X1 i_158 (.A(n_220), .B1(n_217), .B2(n_219), .ZN(n_221));
   NAND2_X1 i_159 (.A1(A[0]), .A2(B[10]), .ZN(n_223));
   XNOR2_X1 i_160 (.A(n_374), .B(n_223), .ZN(n_224));
   XOR2_X1 i_161 (.A(n_224), .B(n_385), .Z(n_225));
   XOR2_X1 i_162 (.A(n_376), .B(n_390), .Z(n_231));
   XOR2_X1 i_163 (.A(n_225), .B(n_231), .Z(n_232));
   AOI22_X1 i_164 (.A1(n_186), .A2(n_190), .B1(n_184), .B2(n_185), .ZN(n_233));
   XNOR2_X1 i_165 (.A(n_232), .B(n_233), .ZN(n_234));
   XOR2_X1 i_166 (.A(n_221), .B(n_234), .Z(n_235));
   INV_X1 i_167 (.A(n_162), .ZN(n_236));
   INV_X1 i_168 (.A(n_193), .ZN(n_237));
   INV_X1 i_169 (.A(n_194), .ZN(n_238));
   AOI21_X1 i_170 (.A(n_237), .B1(n_180), .B2(n_238), .ZN(n_239));
   NAND2_X1 i_171 (.A1(n_236), .A2(n_239), .ZN(n_240));
   OAI21_X1 i_172 (.A(n_240), .B1(n_236), .B2(n_239), .ZN(n_241));
   XOR2_X1 i_173 (.A(n_235), .B(n_241), .Z(n_242));
   OAI21_X1 i_174 (.A(n_196), .B1(n_160), .B2(n_197), .ZN(n_243));
   XNOR2_X1 i_175 (.A(n_242), .B(n_243), .ZN(Out[10]));
   AOI22_X1 i_176 (.A1(n_211), .A2(n_216), .B1(n_210), .B2(n_203), .ZN(n_244));
   OAI33_X1 i_177 (.A1(n_214), .A2(n_99), .A3(n_1955), .B1(n_389), .B2(n_423), 
      .B3(n_169), .ZN(n_247));
   AOI21_X1 i_178 (.A(n_199), .B1(n_201), .B2(n_202), .ZN(n_248));
   XNOR2_X1 i_179 (.A(n_247), .B(n_248), .ZN(n_249));
   OAI22_X1 i_180 (.A1(n_224), .A2(n_385), .B1(n_374), .B2(n_223), .ZN(n_250));
   XNOR2_X1 i_181 (.A(n_249), .B(n_250), .ZN(n_251));
   XOR2_X1 i_182 (.A(n_244), .B(n_251), .Z(n_252));
   INV_X1 i_183 (.A(n_233), .ZN(n_253));
   AOI22_X1 i_184 (.A1(n_232), .A2(n_253), .B1(n_231), .B2(n_225), .ZN(n_254));
   XOR2_X1 i_185 (.A(n_252), .B(n_254), .Z(n_255));
   XNOR2_X1 i_186 (.A(n_439), .B(n_437), .ZN(n_271));
   XNOR2_X1 i_187 (.A(n_375), .B(n_355), .ZN(n_288));
   XNOR2_X1 i_188 (.A(n_271), .B(n_288), .ZN(n_289));
   XNOR2_X1 i_189 (.A(n_255), .B(n_289), .ZN(n_290));
   OAI21_X1 i_190 (.A(n_220), .B1(n_221), .B2(n_234), .ZN(n_291));
   NOR2_X1 i_191 (.A1(n_291), .A2(n_240), .ZN(n_292));
   AOI21_X1 i_192 (.A(n_292), .B1(n_240), .B2(n_291), .ZN(n_293));
   XNOR2_X1 i_193 (.A(n_290), .B(n_293), .ZN(n_294));
   AOI22_X1 i_194 (.A1(n_243), .A2(n_242), .B1(n_235), .B2(n_241), .ZN(n_295));
   XOR2_X1 i_195 (.A(n_294), .B(n_295), .Z(Out[11]));
   AOI22_X1 i_196 (.A1(n_252), .A2(n_254), .B1(n_244), .B2(n_251), .ZN(n_296));
   INV_X1 i_197 (.A(n_248), .ZN(n_297));
   AOI22_X1 i_198 (.A1(n_249), .A2(n_250), .B1(n_247), .B2(n_297), .ZN(n_298));
   INV_X1 i_199 (.A(n_198), .ZN(n_299));
   AOI21_X1 i_200 (.A(n_373), .B1(n_371), .B2(n_299), .ZN(n_300));
   AOI21_X1 i_201 (.A(n_369), .B1(n_359), .B2(n_358), .ZN(n_301));
   XNOR2_X1 i_202 (.A(n_300), .B(n_301), .ZN(n_302));
   XNOR2_X1 i_203 (.A(n_298), .B(n_302), .ZN(n_303));
   XNOR2_X1 i_204 (.A(n_321), .B(n_269), .ZN(n_310));
   XOR2_X1 i_205 (.A(n_207), .B(n_208), .Z(n_315));
   XOR2_X1 i_206 (.A(n_310), .B(n_315), .Z(n_316));
   XNOR2_X1 i_207 (.A(n_303), .B(n_316), .ZN(n_317));
   XOR2_X1 i_208 (.A(n_296), .B(n_317), .Z(n_318));
   XOR2_X1 i_209 (.A(n_427), .B(n_354), .Z(n_322));
   XNOR2_X1 i_210 (.A(n_262), .B(n_263), .ZN(n_329));
   OAI21_X1 i_211 (.A(n_174), .B1(n_168), .B2(n_171), .ZN(n_336));
   XOR2_X1 i_212 (.A(n_329), .B(n_336), .Z(n_337));
   XNOR2_X1 i_213 (.A(n_177), .B(n_178), .ZN(n_341));
   XOR2_X1 i_214 (.A(n_337), .B(n_341), .Z(n_342));
   XNOR2_X1 i_215 (.A(n_322), .B(n_342), .ZN(n_343));
   XOR2_X1 i_216 (.A(n_318), .B(n_343), .Z(n_344));
   OAI22_X1 i_217 (.A1(n_255), .A2(n_289), .B1(n_271), .B2(n_288), .ZN(n_345));
   NAND2_X1 i_218 (.A1(n_345), .A2(n_292), .ZN(n_346));
   OAI21_X1 i_219 (.A(n_346), .B1(n_292), .B2(n_345), .ZN(n_347));
   XNOR2_X1 i_220 (.A(n_344), .B(n_347), .ZN(n_348));
   INV_X1 i_221 (.A(n_295), .ZN(n_349));
   INV_X1 i_222 (.A(n_293), .ZN(n_350));
   AOI22_X1 i_223 (.A1(n_349), .A2(n_294), .B1(n_350), .B2(n_290), .ZN(n_351));
   XOR2_X1 i_224 (.A(n_348), .B(n_351), .Z(Out[12]));
   AOI22_X1 i_225 (.A1(n_322), .A2(n_342), .B1(n_427), .B2(n_354), .ZN(n_352));
   OAI22_X1 i_226 (.A1(n_298), .A2(n_302), .B1(n_300), .B2(n_301), .ZN(n_353));
   XOR2_X1 i_227 (.A(n_189), .B(n_212), .Z(n_360));
   XOR2_X1 i_228 (.A(n_353), .B(n_360), .Z(n_361));
   AOI22_X1 i_229 (.A1(n_337), .A2(n_341), .B1(n_329), .B2(n_336), .ZN(n_362));
   XNOR2_X1 i_230 (.A(n_361), .B(n_362), .ZN(n_363));
   XNOR2_X1 i_231 (.A(n_352), .B(n_363), .ZN(n_364));
   AOI22_X1 i_232 (.A1(n_318), .A2(n_343), .B1(n_296), .B2(n_317), .ZN(n_365));
   XOR2_X1 i_233 (.A(n_364), .B(n_365), .Z(n_366));
   INV_X1 i_234 (.A(n_346), .ZN(n_367));
   XOR2_X1 i_235 (.A(n_312), .B(n_305), .Z(n_383));
   XNOR2_X1 i_236 (.A(n_276), .B(n_275), .ZN(n_401));
   XOR2_X1 i_237 (.A(n_383), .B(n_401), .Z(n_402));
   AOI22_X1 i_238 (.A1(n_303), .A2(n_316), .B1(n_310), .B2(n_315), .ZN(n_403));
   XOR2_X1 i_239 (.A(n_402), .B(n_403), .Z(n_404));
   NAND2_X1 i_240 (.A1(n_367), .A2(n_404), .ZN(n_405));
   OAI21_X1 i_241 (.A(n_405), .B1(n_367), .B2(n_404), .ZN(n_406));
   XNOR2_X1 i_242 (.A(n_366), .B(n_406), .ZN(n_407));
   INV_X1 i_243 (.A(n_347), .ZN(n_408));
   AOI22_X1 i_244 (.A1(n_351), .A2(n_348), .B1(n_408), .B2(n_344), .ZN(n_409));
   XOR2_X1 i_245 (.A(n_407), .B(n_409), .Z(Out[13]));
   INV_X1 i_246 (.A(n_352), .ZN(n_410));
   AOI22_X1 i_247 (.A1(n_365), .A2(n_364), .B1(n_410), .B2(n_363), .ZN(n_411));
   INV_X1 i_248 (.A(n_405), .ZN(n_412));
   NAND2_X1 i_249 (.A1(n_411), .A2(n_412), .ZN(n_413));
   OAI21_X1 i_250 (.A(n_413), .B1(n_411), .B2(n_412), .ZN(n_414));
   AOI22_X1 i_251 (.A1(n_403), .A2(n_402), .B1(n_383), .B2(n_401), .ZN(n_415));
   XOR2_X1 i_252 (.A(n_273), .B(n_268), .Z(n_428));
   XNOR2_X1 i_253 (.A(n_415), .B(n_428), .ZN(n_429));
   AOI22_X1 i_254 (.A1(n_361), .A2(n_362), .B1(n_353), .B2(n_360), .ZN(n_430));
   AOI21_X1 i_255 (.A(n_309), .B1(n_307), .B2(n_306), .ZN(n_431));
   AOI21_X1 i_256 (.A(n_281), .B1(n_283), .B2(n_270), .ZN(n_432));
   XNOR2_X1 i_257 (.A(n_431), .B(n_432), .ZN(n_433));
   INV_X1 i_258 (.A(n_286), .ZN(n_434));
   AOI21_X1 i_259 (.A(n_285), .B1(n_434), .B2(n_284), .ZN(n_435));
   XOR2_X1 i_260 (.A(n_433), .B(n_435), .Z(n_436));
   NOR2_X1 i_261 (.A1(n_520), .A2(n_523), .ZN(n_440));
   XOR2_X1 i_262 (.A(n_440), .B(n_517), .Z(n_443));
   NOR2_X1 i_263 (.A1(n_534), .A2(n_537), .ZN(n_447));
   XNOR2_X1 i_264 (.A(n_447), .B(n_287), .ZN(n_448));
   XOR2_X1 i_265 (.A(n_443), .B(n_448), .Z(n_449));
   XNOR2_X1 i_266 (.A(n_436), .B(n_449), .ZN(n_450));
   NAND2_X1 i_267 (.A1(n_430), .A2(n_450), .ZN(n_451));
   OAI21_X1 i_268 (.A(n_451), .B1(n_430), .B2(n_450), .ZN(n_452));
   XOR2_X1 i_269 (.A(n_492), .B(n_489), .Z(n_456));
   XOR2_X1 i_270 (.A(n_466), .B(n_465), .Z(n_463));
   XOR2_X1 i_271 (.A(n_456), .B(n_463), .Z(n_464));
   XNOR2_X1 i_272 (.A(n_541), .B(n_540), .ZN(n_471));
   NAND2_X1 i_273 (.A1(n_464), .A2(n_471), .ZN(n_472));
   OAI21_X1 i_274 (.A(n_472), .B1(n_464), .B2(n_471), .ZN(n_473));
   XNOR2_X1 i_275 (.A(n_452), .B(n_473), .ZN(n_474));
   XOR2_X1 i_276 (.A(n_429), .B(n_474), .Z(n_475));
   XNOR2_X1 i_277 (.A(n_414), .B(n_475), .ZN(n_476));
   OAI22_X1 i_278 (.A1(n_409), .A2(n_407), .B1(n_366), .B2(n_406), .ZN(n_477));
   XOR2_X1 i_279 (.A(n_476), .B(n_477), .Z(Out[14]));
   INV_X1 i_280 (.A(n_414), .ZN(n_478));
   AOI22_X1 i_281 (.A1(n_477), .A2(n_476), .B1(n_478), .B2(n_475), .ZN(n_479));
   INV_X1 i_282 (.A(n_413), .ZN(n_480));
   INV_X1 i_283 (.A(n_415), .ZN(n_481));
   AOI22_X1 i_284 (.A1(n_474), .A2(n_429), .B1(n_481), .B2(n_428), .ZN(n_482));
   INV_X1 i_285 (.A(n_482), .ZN(n_483));
   NAND2_X1 i_286 (.A1(n_480), .A2(n_483), .ZN(n_484));
   OAI21_X1 i_287 (.A(n_484), .B1(n_480), .B2(n_483), .ZN(n_485));
   OAI21_X1 i_288 (.A(n_451), .B1(n_452), .B2(n_473), .ZN(n_486));
   INV_X1 i_289 (.A(n_578), .ZN(n_490));
   NAND2_X1 i_290 (.A1(n_580), .A2(n_490), .ZN(n_491));
   XOR2_X1 i_291 (.A(n_491), .B(n_579), .Z(n_493));
   NAND2_X1 i_292 (.A1(n_571), .A2(n_568), .ZN(n_497));
   XOR2_X1 i_293 (.A(n_497), .B(n_569), .Z(n_499));
   XOR2_X1 i_294 (.A(n_493), .B(n_499), .Z(n_500));
   NAND2_X1 i_295 (.A1(A[0]), .A2(B[15]), .ZN(n_503));
   XOR2_X1 i_296 (.A(n_502), .B(n_503), .Z(n_504));
   XNOR2_X1 i_297 (.A(n_500), .B(n_504), .ZN(n_505));
   OAI21_X1 i_298 (.A(n_472), .B1(n_463), .B2(n_456), .ZN(n_506));
   XOR2_X1 i_299 (.A(n_505), .B(n_506), .Z(n_507));
   AOI22_X1 i_300 (.A1(n_436), .A2(n_449), .B1(n_448), .B2(n_443), .ZN(n_508));
   XOR2_X1 i_301 (.A(n_507), .B(n_508), .Z(n_509));
   XOR2_X1 i_302 (.A(n_486), .B(n_509), .Z(n_510));
   INV_X1 i_303 (.A(n_304), .ZN(n_511));
   AOI22_X1 i_304 (.A1(n_273), .A2(n_268), .B1(n_511), .B2(n_274), .ZN(n_512));
   INV_X1 i_305 (.A(n_431), .ZN(n_513));
   AOI22_X1 i_306 (.A1(n_433), .A2(n_435), .B1(n_513), .B2(n_432), .ZN(n_514));
   XNOR2_X1 i_307 (.A(n_614), .B(n_615), .ZN(n_518));
   XOR2_X1 i_308 (.A(n_514), .B(n_518), .Z(n_519));
   XNOR2_X1 i_309 (.A(n_565), .B(n_566), .ZN(n_525));
   XNOR2_X1 i_310 (.A(n_519), .B(n_525), .ZN(n_526));
   XNOR2_X1 i_311 (.A(n_512), .B(n_526), .ZN(n_527));
   INV_X1 i_312 (.A(n_222), .ZN(n_528));
   AOI22_X1 i_313 (.A1(n_246), .A2(n_267), .B1(n_528), .B2(n_245), .ZN(n_529));
   XOR2_X1 i_314 (.A(n_524), .B(n_516), .Z(n_538));
   XOR2_X1 i_315 (.A(n_529), .B(n_538), .Z(n_539));
   XOR2_X1 i_316 (.A(n_470), .B(n_462), .Z(n_545));
   XOR2_X1 i_317 (.A(n_539), .B(n_545), .Z(n_546));
   XNOR2_X1 i_318 (.A(n_527), .B(n_546), .ZN(n_547));
   XOR2_X1 i_319 (.A(n_510), .B(n_547), .Z(n_548));
   XNOR2_X1 i_320 (.A(n_485), .B(n_548), .ZN(n_549));
   XOR2_X1 i_321 (.A(n_479), .B(n_549), .Z(Out[15]));
   OAI22_X1 i_322 (.A1(n_479), .A2(n_549), .B1(n_485), .B2(n_548), .ZN(n_550));
   INV_X1 i_323 (.A(n_550), .ZN(n_551));
   INV_X1 i_324 (.A(n_512), .ZN(n_552));
   AOI22_X1 i_325 (.A1(n_527), .A2(n_546), .B1(n_552), .B2(n_526), .ZN(n_553));
   AOI22_X1 i_326 (.A1(n_539), .A2(n_545), .B1(n_529), .B2(n_538), .ZN(n_554));
   XNOR2_X1 i_327 (.A(n_495), .B(n_461), .ZN(n_563));
   XNOR2_X1 i_328 (.A(n_772), .B(n_773), .ZN(n_584));
   XOR2_X1 i_329 (.A(n_563), .B(n_584), .Z(n_585));
   XOR2_X1 i_330 (.A(n_554), .B(n_585), .Z(n_586));
   XOR2_X1 i_331 (.A(n_553), .B(n_586), .Z(n_587));
   AOI22_X1 i_332 (.A1(n_500), .A2(n_504), .B1(n_493), .B2(n_499), .ZN(n_588));
   XOR2_X1 i_333 (.A(n_576), .B(n_581), .Z(n_594));
   XNOR2_X1 i_334 (.A(n_588), .B(n_594), .ZN(n_595));
   AOI22_X1 i_335 (.A1(n_519), .A2(n_525), .B1(n_514), .B2(n_518), .ZN(n_596));
   XOR2_X1 i_336 (.A(n_595), .B(n_596), .Z(n_597));
   XOR2_X1 i_337 (.A(n_781), .B(n_782), .Z(n_617));
   XOR2_X1 i_338 (.A(n_597), .B(n_617), .Z(n_618));
   AOI22_X1 i_339 (.A1(n_507), .A2(n_508), .B1(n_505), .B2(n_506), .ZN(n_619));
   XOR2_X1 i_340 (.A(n_618), .B(n_619), .Z(n_620));
   NAND2_X1 i_341 (.A1(n_587), .A2(n_620), .ZN(n_621));
   OAI21_X1 i_342 (.A(n_621), .B1(n_587), .B2(n_620), .ZN(n_622));
   NAND2_X1 i_343 (.A1(n_551), .A2(n_622), .ZN(n_623));
   OR2_X1 i_344 (.A1(n_551), .A2(n_622), .ZN(n_624));
   NAND2_X1 i_345 (.A1(n_623), .A2(n_624), .ZN(n_625));
   AOI22_X1 i_346 (.A1(n_510), .A2(n_547), .B1(n_486), .B2(n_509), .ZN(n_626));
   INV_X1 i_347 (.A(n_626), .ZN(n_627));
   NOR2_X1 i_348 (.A1(n_484), .A2(n_627), .ZN(n_628));
   AOI21_X1 i_349 (.A(n_628), .B1(n_484), .B2(n_627), .ZN(n_629));
   XNOR2_X1 i_350 (.A(n_625), .B(n_629), .ZN(Out[16]));
   INV_X1 i_351 (.A(n_624), .ZN(n_630));
   OAI21_X1 i_352 (.A(n_623), .B1(n_630), .B2(n_629), .ZN(n_631));
   OAI21_X1 i_353 (.A(n_621), .B1(n_553), .B2(n_586), .ZN(n_632));
   NAND2_X1 i_354 (.A1(n_628), .A2(n_632), .ZN(n_633));
   OAI21_X1 i_355 (.A(n_633), .B1(n_628), .B2(n_632), .ZN(n_634));
   AOI22_X1 i_356 (.A1(n_618), .A2(n_619), .B1(n_597), .B2(n_617), .ZN(n_635));
   INV_X1 i_357 (.A(n_588), .ZN(n_636));
   AOI22_X1 i_358 (.A1(n_595), .A2(n_596), .B1(n_636), .B2(n_594), .ZN(n_637));
   NAND2_X1 i_359 (.A1(B[10]), .A2(A[8]), .ZN(n_638));
   OR3_X1 i_360 (.A1(n_638), .A2(n_556), .A3(n_426), .ZN(n_639));
   OAI22_X1 i_361 (.A1(n_556), .A2(n_2243), .B1(n_458), .B2(n_426), .ZN(n_641));
   NAND2_X1 i_362 (.A1(n_639), .A2(n_641), .ZN(n_642));
   NAND2_X1 i_363 (.A1(A[6]), .A2(B[11]), .ZN(n_643));
   XNOR2_X1 i_364 (.A(n_642), .B(n_643), .ZN(n_644));
   NOR2_X1 i_365 (.A1(n_1955), .A2(n_1339), .ZN(n_646));
   NOR2_X1 i_366 (.A1(n_169), .A2(n_1235), .ZN(n_648));
   NAND2_X1 i_367 (.A1(n_646), .A2(n_648), .ZN(n_649));
   OAI21_X1 i_368 (.A(n_649), .B1(n_646), .B2(n_648), .ZN(n_650));
   NAND2_X1 i_369 (.A1(B[8]), .A2(A[9]), .ZN(n_651));
   XNOR2_X1 i_370 (.A(n_650), .B(n_651), .ZN(n_652));
   XOR2_X1 i_371 (.A(n_644), .B(n_652), .Z(n_653));
   NAND2_X1 i_372 (.A1(A[4]), .A2(B[13]), .ZN(n_654));
   XNOR2_X1 i_373 (.A(n_599), .B(n_654), .ZN(n_655));
   NAND2_X1 i_374 (.A1(A[3]), .A2(B[14]), .ZN(n_656));
   XNOR2_X1 i_375 (.A(n_655), .B(n_656), .ZN(n_657));
   XOR2_X1 i_376 (.A(n_653), .B(n_657), .Z(n_658));
   XOR2_X1 i_377 (.A(n_637), .B(n_658), .Z(n_659));
   XNOR2_X1 i_378 (.A(n_666), .B(n_671), .ZN(n_672));
   XOR2_X1 i_379 (.A(n_659), .B(n_672), .Z(n_673));
   XOR2_X1 i_380 (.A(n_635), .B(n_673), .Z(n_674));
   XOR2_X1 i_381 (.A(n_611), .B(n_460), .Z(n_688));
   XNOR2_X1 i_382 (.A(n_777), .B(n_783), .ZN(n_697));
   XOR2_X1 i_383 (.A(n_688), .B(n_697), .Z(n_698));
   AOI22_X1 i_384 (.A1(n_554), .A2(n_585), .B1(n_563), .B2(n_584), .ZN(n_699));
   XOR2_X1 i_385 (.A(n_698), .B(n_699), .Z(n_700));
   NAND2_X1 i_386 (.A1(n_674), .A2(n_700), .ZN(n_701));
   OAI21_X1 i_387 (.A(n_701), .B1(n_674), .B2(n_700), .ZN(n_702));
   OR2_X1 i_388 (.A1(n_634), .A2(n_702), .ZN(n_703));
   NAND2_X1 i_389 (.A1(n_634), .A2(n_702), .ZN(n_704));
   NAND2_X1 i_390 (.A1(n_703), .A2(n_704), .ZN(n_705));
   XOR2_X1 i_391 (.A(n_631), .B(n_705), .Z(Out[17]));
   INV_X1 i_392 (.A(n_704), .ZN(n_706));
   OAI21_X1 i_393 (.A(n_703), .B1(n_631), .B2(n_706), .ZN(n_707));
   INV_X1 i_394 (.A(n_707), .ZN(n_708));
   NAND2_X1 i_395 (.A1(n_708), .A2(n_633), .ZN(n_709));
   OR2_X1 i_396 (.A1(n_708), .A2(n_633), .ZN(n_710));
   NAND2_X1 i_397 (.A1(n_709), .A2(n_710), .ZN(n_711));
   AOI22_X1 i_398 (.A1(n_698), .A2(n_699), .B1(n_688), .B2(n_697), .ZN(n_712));
   INV_X1 i_399 (.A(n_582), .ZN(n_713));
   INV_X1 i_400 (.A(n_598), .ZN(n_714));
   AOI22_X1 i_401 (.A1(n_713), .A2(n_605), .B1(n_714), .B2(n_604), .ZN(n_715));
   NAND2_X1 i_402 (.A1(A[5]), .A2(B[14]), .ZN(n_716));
   NOR2_X1 i_403 (.A1(n_654), .A2(n_716), .ZN(n_717));
   AOI22_X1 i_404 (.A1(A[4]), .A2(B[14]), .B1(A[5]), .B2(B[13]), .ZN(n_718));
   NOR2_X1 i_405 (.A1(n_717), .A2(n_718), .ZN(n_719));
   NOR2_X1 i_406 (.A1(n_99), .A2(n_560), .ZN(n_720));
   XNOR2_X1 i_407 (.A(n_719), .B(n_720), .ZN(n_721));
   NAND2_X1 i_408 (.A1(A[2]), .A2(B[17]), .ZN(n_722));
   NOR2_X1 i_409 (.A1(n_607), .A2(n_722), .ZN(n_723));
   AOI22_X1 i_410 (.A1(A[1]), .A2(B[17]), .B1(A[2]), .B2(B[16]), .ZN(n_724));
   NOR2_X1 i_411 (.A1(n_723), .A2(n_724), .ZN(n_725));
   NOR2_X1 i_412 (.A1(n_31), .A2(n_1532), .ZN(n_727));
   XNOR2_X1 i_413 (.A(n_725), .B(n_727), .ZN(n_728));
   XOR2_X1 i_414 (.A(n_721), .B(n_728), .Z(n_729));
   XOR2_X1 i_415 (.A(n_715), .B(n_729), .Z(n_730));
   OR3_X1 i_416 (.A1(n_1116), .A2(n_1955), .A3(n_1339), .ZN(n_732));
   OAI22_X1 i_417 (.A1(n_425), .A2(n_1339), .B1(n_1955), .B2(n_1235), .ZN(n_733));
   NAND2_X1 i_418 (.A1(n_732), .A2(n_733), .ZN(n_734));
   NAND2_X1 i_419 (.A1(A[9]), .A2(B[9]), .ZN(n_735));
   XNOR2_X1 i_420 (.A(n_734), .B(n_735), .ZN(n_736));
   NAND2_X1 i_421 (.A1(B[4]), .A2(A[14]), .ZN(n_738));
   XNOR2_X1 i_422 (.A(n_1128), .B(n_738), .ZN(n_739));
   NAND2_X1 i_423 (.A1(B[6]), .A2(A[12]), .ZN(n_740));
   XNOR2_X1 i_424 (.A(n_739), .B(n_740), .ZN(n_741));
   XOR2_X1 i_425 (.A(n_736), .B(n_741), .Z(n_742));
   NAND2_X1 i_426 (.A1(A[7]), .A2(B[11]), .ZN(n_743));
   XNOR2_X1 i_427 (.A(n_638), .B(n_743), .ZN(n_744));
   NAND2_X1 i_428 (.A1(A[6]), .A2(B[12]), .ZN(n_745));
   XNOR2_X1 i_429 (.A(n_744), .B(n_745), .ZN(n_746));
   XOR2_X1 i_430 (.A(n_742), .B(n_746), .Z(n_747));
   NAND2_X1 i_431 (.A1(n_730), .A2(n_747), .ZN(n_748));
   OAI21_X1 i_432 (.A(n_748), .B1(n_730), .B2(n_747), .ZN(n_749));
   AOI22_X1 i_433 (.A1(n_611), .A2(n_459), .B1(n_606), .B2(n_610), .ZN(n_751));
   XOR2_X1 i_434 (.A(n_749), .B(n_751), .Z(n_752));
   XOR2_X1 i_435 (.A(n_712), .B(n_752), .Z(n_753));
   AOI22_X1 i_436 (.A1(n_659), .A2(n_672), .B1(n_637), .B2(n_658), .ZN(n_754));
   OAI21_X1 i_437 (.A(n_639), .B1(n_642), .B2(n_643), .ZN(n_755));
   OAI21_X1 i_438 (.A(n_649), .B1(n_650), .B2(n_651), .ZN(n_756));
   XOR2_X1 i_439 (.A(n_755), .B(n_756), .Z(n_757));
   OAI22_X1 i_440 (.A1(n_655), .A2(n_656), .B1(n_599), .B2(n_654), .ZN(n_758));
   XNOR2_X1 i_441 (.A(n_757), .B(n_758), .ZN(n_759));
   XNOR2_X1 i_442 (.A(n_849), .B(n_848), .ZN(n_764));
   XOR2_X1 i_443 (.A(n_759), .B(n_764), .Z(n_765));
   AOI22_X1 i_444 (.A1(n_653), .A2(n_657), .B1(n_644), .B2(n_652), .ZN(n_766));
   XOR2_X1 i_445 (.A(n_765), .B(n_766), .Z(n_767));
   XOR2_X1 i_446 (.A(n_754), .B(n_767), .Z(n_768));
   XOR2_X1 i_447 (.A(n_802), .B(n_831), .Z(n_785));
   XNOR2_X1 i_448 (.A(n_768), .B(n_785), .ZN(n_786));
   XNOR2_X1 i_449 (.A(n_753), .B(n_786), .ZN(n_787));
   OAI21_X1 i_450 (.A(n_701), .B1(n_635), .B2(n_673), .ZN(n_788));
   XNOR2_X1 i_451 (.A(n_787), .B(n_788), .ZN(n_789));
   XOR2_X1 i_452 (.A(n_711), .B(n_789), .Z(Out[18]));
   NAND2_X1 i_453 (.A1(n_787), .A2(n_788), .ZN(n_790));
   INV_X1 i_454 (.A(n_709), .ZN(n_791));
   OAI211_X1 i_455 (.A(n_710), .B(n_790), .C1(n_791), .C2(n_789), .ZN(n_792));
   INV_X1 i_456 (.A(n_766), .ZN(n_793));
   AOI22_X1 i_457 (.A1(n_765), .A2(n_793), .B1(n_764), .B2(n_759), .ZN(n_794));
   AOI22_X1 i_458 (.A1(n_715), .A2(n_729), .B1(n_721), .B2(n_728), .ZN(n_795));
   XOR2_X1 i_459 (.A(n_794), .B(n_795), .Z(n_796));
   AOI22_X1 i_460 (.A1(n_757), .A2(n_758), .B1(n_756), .B2(n_755), .ZN(n_797));
   AOI21_X1 i_461 (.A(n_717), .B1(n_719), .B2(n_720), .ZN(n_798));
   AOI21_X1 i_462 (.A(n_723), .B1(n_725), .B2(n_727), .ZN(n_799));
   XNOR2_X1 i_463 (.A(n_798), .B(n_799), .ZN(n_800));
   XNOR2_X1 i_464 (.A(n_797), .B(n_800), .ZN(n_801));
   NAND2_X1 i_465 (.A1(A[0]), .A2(B[19]), .ZN(n_803));
   XNOR2_X1 i_466 (.A(n_913), .B(n_803), .ZN(n_804));
   XNOR2_X1 i_467 (.A(n_804), .B(n_722), .ZN(n_805));
   NAND2_X1 i_468 (.A1(A[4]), .A2(B[15]), .ZN(n_806));
   XNOR2_X1 i_469 (.A(n_716), .B(n_806), .ZN(n_807));
   NAND2_X1 i_470 (.A1(A[3]), .A2(B[16]), .ZN(n_808));
   XNOR2_X1 i_471 (.A(n_807), .B(n_808), .ZN(n_809));
   XOR2_X1 i_472 (.A(n_805), .B(n_809), .Z(n_810));
   XOR2_X1 i_473 (.A(n_801), .B(n_810), .Z(n_811));
   XOR2_X1 i_474 (.A(n_796), .B(n_811), .Z(n_812));
   AOI22_X1 i_475 (.A1(n_742), .A2(n_746), .B1(n_736), .B2(n_741), .ZN(n_813));
   OAI21_X1 i_476 (.A(n_732), .B1(n_734), .B2(n_735), .ZN(n_814));
   OAI22_X1 i_477 (.A1(n_739), .A2(n_740), .B1(n_1128), .B2(n_738), .ZN(n_815));
   XOR2_X1 i_478 (.A(n_814), .B(n_815), .Z(n_816));
   OAI33_X1 i_479 (.A1(n_744), .A2(n_170), .A3(n_1676), .B1(n_743), .B2(n_2243), 
      .B3(n_458), .ZN(n_818));
   XOR2_X1 i_480 (.A(n_816), .B(n_818), .Z(n_819));
   XOR2_X1 i_481 (.A(n_813), .B(n_819), .Z(n_820));
   INV_X1 i_482 (.A(n_750), .ZN(n_821));
   OAI22_X1 i_483 (.A1(n_694), .A2(n_761), .B1(n_760), .B2(n_821), .ZN(n_822));
   XNOR2_X1 i_484 (.A(n_820), .B(n_822), .ZN(n_823));
   OR2_X1 i_485 (.A1(n_812), .A2(n_823), .ZN(n_824));
   NAND2_X1 i_486 (.A1(n_812), .A2(n_823), .ZN(n_825));
   NAND2_X1 i_487 (.A1(n_824), .A2(n_825), .ZN(n_826));
   OAI21_X1 i_488 (.A(n_748), .B1(n_751), .B2(n_749), .ZN(n_827));
   XOR2_X1 i_489 (.A(n_826), .B(n_827), .Z(n_828));
   XOR2_X1 i_490 (.A(n_1120), .B(n_1017), .Z(n_854));
   XNOR2_X1 i_491 (.A(n_1115), .B(n_1114), .ZN(n_858));
   XOR2_X1 i_492 (.A(n_854), .B(n_858), .Z(n_859));
   NOR2_X1 i_493 (.A1(n_743), .A2(n_1008), .ZN(n_861));
   AOI22_X1 i_494 (.A1(A[7]), .A2(B[12]), .B1(A[8]), .B2(B[11]), .ZN(n_862));
   NOR2_X1 i_495 (.A1(n_861), .A2(n_862), .ZN(n_863));
   NOR2_X1 i_496 (.A1(n_170), .A2(n_229), .ZN(n_864));
   XNOR2_X1 i_497 (.A(n_863), .B(n_864), .ZN(n_865));
   XOR2_X1 i_498 (.A(n_859), .B(n_865), .Z(n_866));
   NAND2_X1 i_499 (.A1(n_833), .A2(n_866), .ZN(n_867));
   OAI21_X1 i_500 (.A(n_867), .B1(n_866), .B2(n_833), .ZN(n_868));
   XNOR2_X1 i_501 (.A(n_832), .B(n_868), .ZN(n_869));
   XNOR2_X1 i_502 (.A(n_828), .B(n_869), .ZN(n_870));
   AOI22_X1 i_503 (.A1(n_768), .A2(n_785), .B1(n_754), .B2(n_767), .ZN(n_871));
   XOR2_X1 i_504 (.A(n_870), .B(n_871), .Z(n_872));
   AOI22_X1 i_505 (.A1(n_786), .A2(n_753), .B1(n_712), .B2(n_752), .ZN(n_873));
   NAND2_X1 i_506 (.A1(n_872), .A2(n_873), .ZN(n_874));
   OAI21_X1 i_507 (.A(n_874), .B1(n_872), .B2(n_873), .ZN(n_875));
   INV_X1 i_508 (.A(n_875), .ZN(n_876));
   NOR2_X1 i_509 (.A1(n_710), .A2(n_790), .ZN(n_877));
   OAI21_X1 i_510 (.A(n_792), .B1(n_876), .B2(n_877), .ZN(n_878));
   OAI21_X1 i_511 (.A(n_878), .B1(n_792), .B2(n_876), .ZN(n_879));
   INV_X1 i_512 (.A(n_877), .ZN(n_880));
   OAI21_X1 i_513 (.A(n_879), .B1(n_875), .B2(n_880), .ZN(Out[19]));
   AOI22_X1 i_514 (.A1(n_818), .A2(n_816), .B1(n_815), .B2(n_814), .ZN(n_881));
   AOI21_X1 i_515 (.A(n_843), .B1(n_846), .B2(n_844), .ZN(n_882));
   XNOR2_X1 i_516 (.A(n_881), .B(n_882), .ZN(n_883));
   XNOR2_X1 i_517 (.A(n_990), .B(n_989), .ZN(n_890));
   XNOR2_X1 i_518 (.A(n_883), .B(n_890), .ZN(n_891));
   AOI22_X1 i_519 (.A1(n_840), .A2(n_834), .B1(n_847), .B2(n_841), .ZN(n_892));
   AOI22_X1 i_520 (.A1(n_859), .A2(n_865), .B1(n_854), .B2(n_858), .ZN(n_893));
   XNOR2_X1 i_521 (.A(n_892), .B(n_893), .ZN(n_894));
   XNOR2_X1 i_522 (.A(n_891), .B(n_894), .ZN(n_895));
   XOR2_X1 i_523 (.A(n_1013), .B(n_1011), .Z(n_900));
   XNOR2_X1 i_524 (.A(n_995), .B(n_994), .ZN(n_907));
   XOR2_X1 i_525 (.A(n_900), .B(n_907), .Z(n_908));
   XOR2_X1 i_526 (.A(n_1022), .B(n_1021), .Z(n_914));
   XOR2_X1 i_527 (.A(n_908), .B(n_914), .Z(n_915));
   XOR2_X1 i_528 (.A(n_895), .B(n_915), .Z(n_916));
   OAI22_X1 i_529 (.A1(n_797), .A2(n_800), .B1(n_798), .B2(n_799), .ZN(n_917));
   OAI22_X1 i_530 (.A1(n_804), .A2(n_722), .B1(n_913), .B2(n_803), .ZN(n_918));
   AOI21_X1 i_531 (.A(n_861), .B1(n_863), .B2(n_864), .ZN(n_919));
   XNOR2_X1 i_532 (.A(n_918), .B(n_919), .ZN(n_920));
   OAI22_X1 i_533 (.A1(n_807), .A2(n_808), .B1(n_716), .B2(n_806), .ZN(n_921));
   XOR2_X1 i_534 (.A(n_920), .B(n_921), .Z(n_922));
   XOR2_X1 i_535 (.A(n_917), .B(n_922), .Z(n_923));
   XOR2_X1 i_536 (.A(n_1117), .B(n_1113), .Z(n_930));
   XNOR2_X1 i_537 (.A(n_923), .B(n_930), .ZN(n_931));
   XNOR2_X1 i_538 (.A(n_916), .B(n_931), .ZN(n_932));
   INV_X1 i_539 (.A(n_825), .ZN(n_933));
   OAI21_X1 i_540 (.A(n_824), .B1(n_933), .B2(n_827), .ZN(n_934));
   NAND2_X1 i_541 (.A1(n_932), .A2(n_934), .ZN(n_935));
   OAI21_X1 i_542 (.A(n_935), .B1(n_932), .B2(n_934), .ZN(n_936));
   AOI22_X1 i_543 (.A1(n_820), .A2(n_822), .B1(n_819), .B2(n_813), .ZN(n_937));
   XNOR2_X1 i_544 (.A(n_924), .B(n_906), .ZN(n_956));
   XNOR2_X1 i_545 (.A(n_937), .B(n_956), .ZN(n_957));
   AOI22_X1 i_546 (.A1(n_801), .A2(n_810), .B1(n_809), .B2(n_805), .ZN(n_958));
   XOR2_X1 i_547 (.A(n_957), .B(n_958), .Z(n_959));
   OAI21_X1 i_548 (.A(n_867), .B1(n_832), .B2(n_868), .ZN(n_960));
   INV_X1 i_549 (.A(n_794), .ZN(n_961));
   INV_X1 i_550 (.A(n_795), .ZN(n_962));
   AOI22_X1 i_551 (.A1(n_796), .A2(n_811), .B1(n_961), .B2(n_962), .ZN(n_963));
   XOR2_X1 i_552 (.A(n_960), .B(n_963), .Z(n_964));
   XOR2_X1 i_553 (.A(n_959), .B(n_964), .Z(n_965));
   XNOR2_X1 i_554 (.A(n_936), .B(n_965), .ZN(n_966));
   NOR2_X1 i_555 (.A1(n_878), .A2(n_966), .ZN(n_967));
   INV_X1 i_556 (.A(n_967), .ZN(n_968));
   NAND2_X1 i_557 (.A1(n_878), .A2(n_966), .ZN(n_969));
   NAND2_X1 i_558 (.A1(n_968), .A2(n_969), .ZN(n_970));
   INV_X1 i_559 (.A(n_871), .ZN(n_971));
   OAI22_X1 i_560 (.A1(n_870), .A2(n_971), .B1(n_828), .B2(n_869), .ZN(n_972));
   NOR2_X1 i_561 (.A1(n_874), .A2(n_972), .ZN(n_973));
   AOI21_X1 i_562 (.A(n_973), .B1(n_874), .B2(n_972), .ZN(n_974));
   XNOR2_X1 i_563 (.A(n_970), .B(n_974), .ZN(Out[20]));
   AOI21_X1 i_564 (.A(n_967), .B1(n_974), .B2(n_969), .ZN(n_975));
   INV_X1 i_565 (.A(n_912), .ZN(n_976));
   NAND2_X1 i_566 (.A1(n_909), .A2(n_976), .ZN(n_977));
   OAI33_X1 i_567 (.A1(n_928), .A2(n_99), .A3(n_1232), .B1(n_939), .B2(n_423), 
      .B3(n_560), .ZN(n_979));
   XOR2_X1 i_568 (.A(n_977), .B(n_979), .Z(n_980));
   INV_X1 i_569 (.A(n_919), .ZN(n_981));
   AOI22_X1 i_570 (.A1(n_920), .A2(n_921), .B1(n_918), .B2(n_981), .ZN(n_982));
   XNOR2_X1 i_571 (.A(n_980), .B(n_982), .ZN(n_983));
   XNOR2_X1 i_572 (.A(n_983), .B(n_901), .ZN(n_997));
   INV_X1 i_573 (.A(n_1052), .ZN(n_1010));
   NAND2_X1 i_574 (.A1(n_1010), .A2(n_1053), .ZN(n_1012));
   XOR2_X1 i_575 (.A(n_1012), .B(n_1035), .Z(n_1019));
   XOR2_X1 i_576 (.A(n_997), .B(n_1019), .Z(n_1020));
   XNOR2_X1 i_577 (.A(n_1103), .B(n_1097), .ZN(n_1037));
   XNOR2_X1 i_578 (.A(n_1020), .B(n_1037), .ZN(n_1038));
   INV_X1 i_579 (.A(n_937), .ZN(n_1039));
   AOI22_X1 i_580 (.A1(n_957), .A2(n_958), .B1(n_1039), .B2(n_956), .ZN(n_1040));
   XNOR2_X1 i_581 (.A(n_1038), .B(n_1040), .ZN(n_1041));
   AOI22_X1 i_582 (.A1(n_916), .A2(n_931), .B1(n_895), .B2(n_915), .ZN(n_1042));
   XNOR2_X1 i_583 (.A(n_1041), .B(n_1042), .ZN(n_1043));
   INV_X1 i_584 (.A(n_960), .ZN(n_1044));
   OAI22_X1 i_585 (.A1(n_959), .A2(n_964), .B1(n_1044), .B2(n_963), .ZN(n_1045));
   INV_X1 i_586 (.A(n_892), .ZN(n_1046));
   AOI22_X1 i_587 (.A1(n_891), .A2(n_894), .B1(n_1046), .B2(n_893), .ZN(n_1047));
   XNOR2_X1 i_588 (.A(n_940), .B(n_905), .ZN(n_1066));
   XOR2_X1 i_589 (.A(n_1047), .B(n_1066), .Z(n_1067));
   INV_X1 i_590 (.A(n_882), .ZN(n_1068));
   AOI22_X1 i_591 (.A1(n_883), .A2(n_890), .B1(n_881), .B2(n_1068), .ZN(n_1069));
   AOI22_X1 i_592 (.A1(n_908), .A2(n_914), .B1(n_907), .B2(n_900), .ZN(n_1070));
   NAND2_X1 i_593 (.A1(n_1069), .A2(n_1070), .ZN(n_1071));
   OAI21_X1 i_594 (.A(n_1071), .B1(n_1069), .B2(n_1070), .ZN(n_1072));
   AOI22_X1 i_595 (.A1(n_923), .A2(n_930), .B1(n_917), .B2(n_922), .ZN(n_1073));
   XNOR2_X1 i_596 (.A(n_1072), .B(n_1073), .ZN(n_1074));
   XOR2_X1 i_597 (.A(n_1067), .B(n_1074), .Z(n_1075));
   XNOR2_X1 i_598 (.A(n_1045), .B(n_1075), .ZN(n_1076));
   XOR2_X1 i_599 (.A(n_1043), .B(n_1076), .Z(n_1077));
   OAI21_X1 i_600 (.A(n_935), .B1(n_936), .B2(n_965), .ZN(n_1078));
   NAND2_X1 i_601 (.A1(n_1077), .A2(n_1078), .ZN(n_1079));
   OAI21_X1 i_602 (.A(n_1079), .B1(n_1077), .B2(n_1078), .ZN(n_1080));
   INV_X1 i_603 (.A(n_973), .ZN(n_1081));
   AND2_X1 i_604 (.A1(n_1080), .A2(n_1081), .ZN(n_1082));
   NOR2_X1 i_605 (.A1(n_1080), .A2(n_1081), .ZN(n_1083));
   NOR2_X1 i_606 (.A1(n_1082), .A2(n_1083), .ZN(n_1084));
   XNOR2_X1 i_607 (.A(n_975), .B(n_1084), .ZN(Out[21]));
   INV_X1 i_608 (.A(n_1083), .ZN(n_1085));
   OAI21_X1 i_609 (.A(n_1085), .B1(n_975), .B2(n_1082), .ZN(n_1086));
   INV_X1 i_610 (.A(n_1079), .ZN(n_1087));
   NOR2_X1 i_611 (.A1(n_1086), .A2(n_1087), .ZN(n_1088));
   INV_X1 i_612 (.A(n_1088), .ZN(n_1089));
   NAND2_X1 i_613 (.A1(n_1086), .A2(n_1087), .ZN(n_1090));
   NAND2_X1 i_614 (.A1(n_1089), .A2(n_1090), .ZN(n_1091));
   INV_X1 i_615 (.A(n_1040), .ZN(n_1092));
   AOI22_X1 i_616 (.A1(n_1041), .A2(n_1042), .B1(n_1038), .B2(n_1092), .ZN(
      n_1093));
   AOI22_X1 i_617 (.A1(n_1020), .A2(n_1037), .B1(n_997), .B2(n_1019), .ZN(n_1094));
   XNOR2_X1 i_618 (.A(n_1032), .B(n_1096), .ZN(n_1105));
   OAI21_X1 i_619 (.A(n_1071), .B1(n_1072), .B2(n_1073), .ZN(n_1106));
   XOR2_X1 i_620 (.A(n_1105), .B(n_1106), .Z(n_1107));
   XNOR2_X1 i_621 (.A(n_1094), .B(n_1107), .ZN(n_1108));
   XOR2_X1 i_622 (.A(n_1093), .B(n_1108), .Z(n_1109));
   AOI22_X1 i_623 (.A1(n_983), .A2(n_901), .B1(n_887), .B2(n_899), .ZN(n_1123));
   XNOR2_X1 i_624 (.A(n_903), .B(n_1123), .ZN(n_1124));
   INV_X1 i_625 (.A(n_982), .ZN(n_1125));
   AOI22_X1 i_626 (.A1(n_980), .A2(n_1125), .B1(n_979), .B2(n_977), .ZN(n_1126));
   NAND2_X1 i_627 (.A1(A[0]), .A2(B[22]), .ZN(n_1127));
   NAND3_X1 i_628 (.A1(n_1530), .A2(A[1]), .A3(B[20]), .ZN(n_1130));
   INV_X1 i_629 (.A(n_1130), .ZN(n_1131));
   AOI22_X1 i_630 (.A1(A[1]), .A2(B[21]), .B1(A[2]), .B2(B[20]), .ZN(n_1132));
   OAI21_X1 i_631 (.A(n_1127), .B1(n_1131), .B2(n_1132), .ZN(n_1133));
   OR3_X1 i_632 (.A1(n_1131), .A2(n_1132), .A3(n_1127), .ZN(n_1134));
   NAND2_X1 i_633 (.A1(n_1133), .A2(n_1134), .ZN(n_1135));
   XOR2_X1 i_634 (.A(n_1126), .B(n_1135), .Z(n_1136));
   AOI21_X1 i_635 (.A(n_1050), .B1(n_1048), .B2(n_1036), .ZN(n_1137));
   AOI21_X1 i_636 (.A(n_884), .B1(n_860), .B2(n_855), .ZN(n_1138));
   XNOR2_X1 i_637 (.A(n_1137), .B(n_1138), .ZN(n_1139));
   AOI21_X1 i_638 (.A(n_896), .B1(n_902), .B2(n_888), .ZN(n_1140));
   XNOR2_X1 i_639 (.A(n_1139), .B(n_1140), .ZN(n_1141));
   XOR2_X1 i_640 (.A(n_1136), .B(n_1141), .Z(n_1142));
   XNOR2_X1 i_641 (.A(n_1301), .B(n_1300), .ZN(n_1149));
   XNOR2_X1 i_642 (.A(n_1296), .B(n_1295), .ZN(n_1155));
   XOR2_X1 i_643 (.A(n_1149), .B(n_1155), .Z(n_1156));
   XOR2_X1 i_644 (.A(n_1289), .B(n_1173), .Z(n_1162));
   XOR2_X1 i_645 (.A(n_1156), .B(n_1162), .Z(n_1163));
   XNOR2_X1 i_646 (.A(n_1051), .B(n_1231), .ZN(n_1165));
   NAND2_X1 i_647 (.A1(A[6]), .A2(B[16]), .ZN(n_1166));
   XNOR2_X1 i_648 (.A(n_1165), .B(n_1166), .ZN(n_1167));
   NAND2_X1 i_649 (.A1(B[11]), .A2(A[11]), .ZN(n_1168));
   XNOR2_X1 i_650 (.A(n_1060), .B(n_1168), .ZN(n_1169));
   NAND2_X1 i_651 (.A1(A[9]), .A2(B[13]), .ZN(n_1170));
   XNOR2_X1 i_652 (.A(n_1169), .B(n_1170), .ZN(n_1171));
   XOR2_X1 i_653 (.A(n_1167), .B(n_1171), .Z(n_1172));
   XNOR2_X1 i_654 (.A(n_889), .B(n_1209), .ZN(n_1174));
   NAND2_X1 i_655 (.A1(A[3]), .A2(B[19]), .ZN(n_1175));
   XNOR2_X1 i_656 (.A(n_1174), .B(n_1175), .ZN(n_1176));
   XOR2_X1 i_657 (.A(n_1172), .B(n_1176), .Z(n_1177));
   XOR2_X1 i_658 (.A(n_1163), .B(n_1177), .Z(n_1178));
   XNOR2_X1 i_659 (.A(n_1142), .B(n_1178), .ZN(n_1179));
   XOR2_X1 i_660 (.A(n_1124), .B(n_1179), .Z(n_1180));
   AOI22_X1 i_661 (.A1(n_1067), .A2(n_1074), .B1(n_1047), .B2(n_1066), .ZN(
      n_1181));
   XNOR2_X1 i_662 (.A(n_1180), .B(n_1181), .ZN(n_1182));
   XNOR2_X1 i_663 (.A(n_1109), .B(n_1182), .ZN(n_1183));
   OAI22_X1 i_664 (.A1(n_1043), .A2(n_1076), .B1(n_1045), .B2(n_1075), .ZN(
      n_1184));
   NAND2_X1 i_665 (.A1(n_1183), .A2(n_1184), .ZN(n_1185));
   OAI21_X1 i_666 (.A(n_1185), .B1(n_1184), .B2(n_1183), .ZN(n_1186));
   XOR2_X1 i_667 (.A(n_1091), .B(n_1186), .Z(Out[22]));
   OAI21_X1 i_668 (.A(n_1090), .B1(n_1088), .B2(n_1186), .ZN(n_1187));
   AOI22_X1 i_669 (.A1(n_1109), .A2(n_1182), .B1(n_1093), .B2(n_1108), .ZN(
      n_1188));
   AOI22_X1 i_670 (.A1(n_1136), .A2(n_1141), .B1(n_1126), .B2(n_1135), .ZN(
      n_1189));
   XNOR2_X1 i_671 (.A(n_1200), .B(n_1199), .ZN(n_1195));
   XNOR2_X1 i_672 (.A(n_1226), .B(n_1225), .ZN(n_1201));
   XOR2_X1 i_673 (.A(n_1195), .B(n_1201), .Z(n_1202));
   XNOR2_X1 i_674 (.A(n_1260), .B(n_1259), .ZN(n_1206));
   XOR2_X1 i_675 (.A(n_1202), .B(n_1206), .Z(n_1207));
   XNOR2_X1 i_676 (.A(n_1189), .B(n_1207), .ZN(n_1208));
   XOR2_X1 i_677 (.A(n_1208), .B(n_1031), .Z(n_1210));
   AOI22_X1 i_678 (.A1(n_903), .A2(n_1123), .B1(n_904), .B2(n_944), .ZN(n_1211));
   NOR2_X1 i_679 (.A1(n_1329), .A2(n_1327), .ZN(n_1215));
   XOR2_X1 i_680 (.A(n_1215), .B(n_949), .Z(n_1216));
   INV_X1 i_681 (.A(n_948), .ZN(n_1217));
   AOI21_X1 i_682 (.A(n_947), .B1(n_950), .B2(n_1217), .ZN(n_1218));
   XOR2_X1 i_683 (.A(n_1216), .B(n_1218), .Z(n_1219));
   XNOR2_X1 i_684 (.A(n_1192), .B(n_1191), .ZN(n_1223));
   XOR2_X1 i_685 (.A(n_1219), .B(n_1223), .Z(n_1224));
   XOR2_X1 i_686 (.A(n_1158), .B(n_1157), .Z(n_1229));
   XNOR2_X1 i_687 (.A(n_1150), .B(n_1148), .ZN(n_1233));
   XOR2_X1 i_688 (.A(n_1229), .B(n_1233), .Z(n_1234));
   INV_X1 i_689 (.A(n_1221), .ZN(n_1237));
   NAND2_X1 i_690 (.A1(n_1220), .A2(n_1237), .ZN(n_1238));
   XNOR2_X1 i_691 (.A(n_1238), .B(n_1214), .ZN(n_1240));
   XNOR2_X1 i_692 (.A(n_1234), .B(n_1240), .ZN(n_1241));
   XOR2_X1 i_693 (.A(n_1224), .B(n_1241), .Z(n_1242));
   XOR2_X1 i_694 (.A(n_1211), .B(n_1242), .Z(n_1243));
   XOR2_X1 i_695 (.A(n_1210), .B(n_1243), .Z(n_1244));
   AOI22_X1 i_696 (.A1(n_1094), .A2(n_1107), .B1(n_1106), .B2(n_1105), .ZN(
      n_1245));
   XOR2_X1 i_697 (.A(n_1244), .B(n_1245), .Z(n_1246));
   AOI22_X1 i_698 (.A1(n_1180), .A2(n_1181), .B1(n_1179), .B2(n_1124), .ZN(
      n_1247));
   AOI22_X1 i_699 (.A1(n_1156), .A2(n_1162), .B1(n_1149), .B2(n_1155), .ZN(
      n_1248));
   INV_X1 i_700 (.A(n_999), .ZN(n_1249));
   AOI22_X1 i_701 (.A1(n_955), .A2(n_945), .B1(n_1249), .B2(n_978), .ZN(n_1250));
   XNOR2_X1 i_702 (.A(n_1248), .B(n_1250), .ZN(n_1251));
   INV_X1 i_703 (.A(n_1137), .ZN(n_1252));
   AOI22_X1 i_704 (.A1(n_1139), .A2(n_1140), .B1(n_1252), .B2(n_1138), .ZN(
      n_1253));
   AND2_X1 i_705 (.A1(n_1134), .A2(n_1130), .ZN(n_1254));
   XOR2_X1 i_706 (.A(n_1253), .B(n_1254), .Z(n_1255));
   AOI22_X1 i_707 (.A1(n_1061), .A2(n_1056), .B1(n_1063), .B2(n_1062), .ZN(
      n_1256));
   XNOR2_X1 i_708 (.A(n_1255), .B(n_1256), .ZN(n_1257));
   XOR2_X1 i_709 (.A(n_1251), .B(n_1257), .Z(n_1258));
   XOR2_X1 i_710 (.A(n_1292), .B(n_1264), .Z(n_1265));
   OAI33_X1 i_711 (.A1(n_1174), .A2(n_99), .A3(n_1711), .B1(n_1209), .B2(n_423), 
      .B3(n_1232), .ZN(n_1267));
   OAI22_X1 i_712 (.A1(n_1169), .A2(n_1170), .B1(n_1060), .B2(n_1168), .ZN(
      n_1268));
   OAI22_X1 i_713 (.A1(n_1165), .A2(n_1166), .B1(n_1051), .B2(n_1231), .ZN(
      n_1269));
   XOR2_X1 i_714 (.A(n_1268), .B(n_1269), .Z(n_1270));
   XNOR2_X1 i_715 (.A(n_1267), .B(n_1270), .ZN(n_1271));
   XOR2_X1 i_716 (.A(n_1265), .B(n_1271), .Z(n_1272));
   AOI22_X1 i_717 (.A1(n_1172), .A2(n_1176), .B1(n_1171), .B2(n_1167), .ZN(
      n_1273));
   XOR2_X1 i_718 (.A(n_1272), .B(n_1273), .Z(n_1274));
   XOR2_X1 i_719 (.A(n_1258), .B(n_1274), .Z(n_1275));
   AOI22_X1 i_720 (.A1(n_1142), .A2(n_1178), .B1(n_1163), .B2(n_1177), .ZN(
      n_1276));
   XNOR2_X1 i_721 (.A(n_1275), .B(n_1276), .ZN(n_1277));
   XOR2_X1 i_722 (.A(n_1247), .B(n_1277), .Z(n_1278));
   XOR2_X1 i_723 (.A(n_1246), .B(n_1278), .Z(n_1279));
   XNOR2_X1 i_724 (.A(n_1188), .B(n_1279), .ZN(n_1280));
   XOR2_X1 i_725 (.A(n_1280), .B(n_1185), .Z(n_1281));
   XNOR2_X1 i_726 (.A(n_1187), .B(n_1281), .ZN(Out[23]));
   OAI21_X1 i_727 (.A(n_1280), .B1(n_1187), .B2(n_1281), .ZN(n_1282));
   INV_X1 i_728 (.A(n_1188), .ZN(n_1283));
   OAI21_X1 i_729 (.A(n_1282), .B1(n_1283), .B2(n_1279), .ZN(n_1284));
   NOR4_X1 i_730 (.A1(n_1090), .A2(n_1185), .A3(n_1283), .A4(n_1279), .ZN(n_1285));
   INV_X1 i_731 (.A(n_1285), .ZN(n_1286));
   NAND2_X1 i_732 (.A1(n_1284), .A2(n_1286), .ZN(n_1287));
   AOI22_X1 i_733 (.A1(n_1202), .A2(n_1206), .B1(n_1201), .B2(n_1195), .ZN(
      n_1288));
   XOR2_X1 i_734 (.A(n_1288), .B(n_1144), .Z(n_1304));
   INV_X1 i_735 (.A(n_1189), .ZN(n_1306));
   AOI22_X1 i_736 (.A1(n_1208), .A2(n_1030), .B1(n_1306), .B2(n_1207), .ZN(
      n_1307));
   XOR2_X1 i_737 (.A(n_1304), .B(n_1307), .Z(n_1308));
   AOI22_X1 i_738 (.A1(n_1211), .A2(n_1242), .B1(n_1241), .B2(n_1224), .ZN(
      n_1309));
   XOR2_X1 i_739 (.A(n_1308), .B(n_1309), .Z(n_1310));
   INV_X1 i_740 (.A(n_1245), .ZN(n_1311));
   AOI22_X1 i_741 (.A1(n_1244), .A2(n_1311), .B1(n_1210), .B2(n_1243), .ZN(
      n_1312));
   XOR2_X1 i_742 (.A(n_1310), .B(n_1312), .Z(n_1313));
   AOI22_X1 i_743 (.A1(n_1276), .A2(n_1275), .B1(n_1258), .B2(n_1274), .ZN(
      n_1314));
   INV_X1 i_744 (.A(n_1273), .ZN(n_1315));
   AOI22_X1 i_745 (.A1(n_1272), .A2(n_1315), .B1(n_1271), .B2(n_1265), .ZN(
      n_1316));
   XOR2_X1 i_746 (.A(n_1418), .B(n_1420), .Z(n_1335));
   XOR2_X1 i_747 (.A(n_1316), .B(n_1335), .Z(n_1336));
   AOI22_X1 i_748 (.A1(n_1255), .A2(n_1256), .B1(n_1253), .B2(n_1254), .ZN(
      n_1337));
   NAND2_X1 i_749 (.A1(n_1479), .A2(n_1481), .ZN(n_1340));
   XNOR2_X1 i_750 (.A(n_1340), .B(n_1478), .ZN(n_1342));
   NAND2_X1 i_751 (.A1(n_1484), .A2(n_1485), .ZN(n_1347));
   XNOR2_X1 i_752 (.A(n_1347), .B(n_1482), .ZN(n_1350));
   XOR2_X1 i_753 (.A(n_1342), .B(n_1350), .Z(n_1351));
   XOR2_X1 i_754 (.A(n_1337), .B(n_1351), .Z(n_1352));
   XOR2_X1 i_755 (.A(n_1336), .B(n_1352), .Z(n_1353));
   XNOR2_X1 i_756 (.A(n_1314), .B(n_1353), .ZN(n_1354));
   INV_X1 i_757 (.A(n_1250), .ZN(n_1355));
   AOI22_X1 i_758 (.A1(n_1251), .A2(n_1257), .B1(n_1355), .B2(n_1248), .ZN(
      n_1356));
   OAI21_X1 i_759 (.A(n_1441), .B1(n_1426), .B2(n_1436), .ZN(n_1379));
   XNOR2_X1 i_760 (.A(n_1356), .B(n_1379), .ZN(n_1380));
   AOI22_X1 i_761 (.A1(n_1270), .A2(n_1267), .B1(n_1268), .B2(n_1269), .ZN(
      n_1385));
   XNOR2_X1 i_762 (.A(n_1236), .B(n_1385), .ZN(n_1386));
   INV_X1 i_763 (.A(n_1218), .ZN(n_1387));
   OAI22_X1 i_764 (.A1(n_1219), .A2(n_1223), .B1(n_1216), .B2(n_1387), .ZN(
      n_1388));
   AOI22_X1 i_765 (.A1(n_1234), .A2(n_1240), .B1(n_1229), .B2(n_1233), .ZN(
      n_1389));
   XOR2_X1 i_766 (.A(n_1388), .B(n_1389), .Z(n_1390));
   XOR2_X1 i_767 (.A(n_1386), .B(n_1390), .Z(n_1391));
   XOR2_X1 i_768 (.A(n_1380), .B(n_1391), .Z(n_1392));
   XNOR2_X1 i_769 (.A(n_1354), .B(n_1392), .ZN(n_1393));
   XOR2_X1 i_770 (.A(n_1313), .B(n_1393), .Z(n_1394));
   AOI22_X1 i_771 (.A1(n_1278), .A2(n_1246), .B1(n_1247), .B2(n_1277), .ZN(
      n_1395));
   INV_X1 i_772 (.A(n_1395), .ZN(n_1396));
   NOR2_X1 i_773 (.A1(n_1394), .A2(n_1396), .ZN(n_1397));
   AOI21_X1 i_774 (.A(n_1397), .B1(n_1396), .B2(n_1394), .ZN(n_1398));
   XNOR2_X1 i_775 (.A(n_1287), .B(n_1398), .ZN(Out[24]));
   OAI21_X1 i_776 (.A(n_1284), .B1(n_1398), .B2(n_1285), .ZN(n_1399));
   INV_X1 i_777 (.A(n_1239), .ZN(n_1400));
   AOI22_X1 i_778 (.A1(n_1236), .A2(n_1385), .B1(n_1263), .B2(n_1400), .ZN(
      n_1401));
   XNOR2_X1 i_779 (.A(n_1362), .B(n_1365), .ZN(n_1407));
   XNOR2_X1 i_780 (.A(n_1401), .B(n_1407), .ZN(n_1408));
   XNOR2_X1 i_781 (.A(n_1501), .B(n_1461), .ZN(n_1416));
   XOR2_X1 i_782 (.A(n_1408), .B(n_1416), .Z(n_1417));
   XOR2_X1 i_783 (.A(n_1423), .B(n_1442), .Z(n_1427));
   XOR2_X1 i_784 (.A(n_1417), .B(n_1427), .Z(n_1428));
   AOI22_X1 i_785 (.A1(n_1336), .A2(n_1352), .B1(n_1316), .B2(n_1335), .ZN(
      n_1429));
   XOR2_X1 i_786 (.A(n_1428), .B(n_1429), .Z(n_1430));
   AOI22_X1 i_787 (.A1(n_1386), .A2(n_1390), .B1(n_1389), .B2(n_1388), .ZN(
      n_1431));
   NAND2_X1 i_788 (.A1(B[6]), .A2(A[19]), .ZN(n_1432));
   XNOR2_X1 i_789 (.A(n_1375), .B(n_1432), .ZN(n_1433));
   NAND2_X1 i_790 (.A1(B[8]), .A2(A[17]), .ZN(n_1434));
   XOR2_X1 i_791 (.A(n_1433), .B(n_1434), .Z(n_1435));
   XNOR2_X1 i_792 (.A(n_1344), .B(n_1631), .ZN(n_1437));
   NAND2_X1 i_793 (.A1(B[11]), .A2(A[14]), .ZN(n_1438));
   XOR2_X1 i_794 (.A(n_1437), .B(n_1438), .Z(n_1439));
   XNOR2_X1 i_795 (.A(n_1435), .B(n_1439), .ZN(n_1440));
   XOR2_X1 i_796 (.A(n_1526), .B(n_1341), .Z(n_1445));
   XNOR2_X1 i_797 (.A(n_1440), .B(n_1445), .ZN(n_1446));
   XNOR2_X1 i_798 (.A(n_1371), .B(n_1372), .ZN(n_1451));
   XNOR2_X1 i_799 (.A(n_1505), .B(n_1504), .ZN(n_1457));
   XOR2_X1 i_800 (.A(n_1451), .B(n_1457), .Z(n_1458));
   NAND2_X1 i_801 (.A1(A[8]), .A2(B[17]), .ZN(n_1462));
   XNOR2_X1 i_802 (.A(n_1522), .B(n_1462), .ZN(n_1463));
   XNOR2_X1 i_803 (.A(n_1458), .B(n_1463), .ZN(n_1464));
   XOR2_X1 i_804 (.A(n_1446), .B(n_1464), .Z(n_1465));
   NAND2_X1 i_805 (.A1(n_1431), .A2(n_1465), .ZN(n_1466));
   OAI21_X1 i_806 (.A(n_1466), .B1(n_1431), .B2(n_1465), .ZN(n_1467));
   XOR2_X1 i_807 (.A(n_1430), .B(n_1467), .Z(n_1468));
   INV_X1 i_808 (.A(n_1314), .ZN(n_1469));
   AOI22_X1 i_809 (.A1(n_1354), .A2(n_1392), .B1(n_1469), .B2(n_1353), .ZN(
      n_1470));
   XNOR2_X1 i_810 (.A(n_1468), .B(n_1470), .ZN(n_1471));
   INV_X1 i_811 (.A(n_1356), .ZN(n_1472));
   AOI22_X1 i_812 (.A1(n_1380), .A2(n_1391), .B1(n_1472), .B2(n_1379), .ZN(
      n_1473));
   INV_X1 i_813 (.A(n_1288), .ZN(n_1474));
   AOI22_X1 i_814 (.A1(n_1144), .A2(n_1474), .B1(n_1196), .B2(n_1145), .ZN(
      n_1475));
   XNOR2_X1 i_815 (.A(n_1326), .B(n_1338), .ZN(n_1486));
   XNOR2_X1 i_816 (.A(n_1475), .B(n_1486), .ZN(n_1487));
   AOI22_X1 i_817 (.A1(n_1337), .A2(n_1351), .B1(n_1350), .B2(n_1342), .ZN(
      n_1488));
   XNOR2_X1 i_818 (.A(n_1487), .B(n_1488), .ZN(n_1489));
   XNOR2_X1 i_819 (.A(n_1473), .B(n_1489), .ZN(n_1490));
   INV_X1 i_820 (.A(n_1309), .ZN(n_1491));
   AOI22_X1 i_821 (.A1(n_1308), .A2(n_1491), .B1(n_1307), .B2(n_1304), .ZN(
      n_1492));
   XOR2_X1 i_822 (.A(n_1490), .B(n_1492), .Z(n_1493));
   XOR2_X1 i_823 (.A(n_1471), .B(n_1493), .Z(n_1494));
   AOI22_X1 i_824 (.A1(n_1313), .A2(n_1393), .B1(n_1312), .B2(n_1310), .ZN(
      n_1495));
   XNOR2_X1 i_825 (.A(n_1494), .B(n_1495), .ZN(n_1496));
   XNOR2_X1 i_826 (.A(n_1496), .B(n_1397), .ZN(n_1497));
   XNOR2_X1 i_827 (.A(n_1399), .B(n_1497), .ZN(Out[25]));
   AOI21_X1 i_828 (.A(n_1496), .B1(n_1399), .B2(n_1497), .ZN(n_1498));
   INV_X1 i_829 (.A(n_1495), .ZN(n_1499));
   AOI22_X1 i_830 (.A1(n_1494), .A2(n_1499), .B1(n_1471), .B2(n_1493), .ZN(
      n_1500));
   XNOR2_X1 i_831 (.A(n_1413), .B(n_1443), .ZN(n_1510));
   OAI21_X1 i_832 (.A(n_1466), .B1(n_1446), .B2(n_1464), .ZN(n_1511));
   XOR2_X1 i_833 (.A(n_1510), .B(n_1511), .Z(n_1512));
   AOI22_X1 i_834 (.A1(n_1428), .A2(n_1429), .B1(n_1417), .B2(n_1427), .ZN(
      n_1513));
   XOR2_X1 i_835 (.A(n_1512), .B(n_1513), .Z(n_1514));
   INV_X1 i_836 (.A(n_1467), .ZN(n_1515));
   OAI22_X1 i_837 (.A1(n_1468), .A2(n_1470), .B1(n_1430), .B2(n_1515), .ZN(
      n_1516));
   XOR2_X1 i_838 (.A(n_1514), .B(n_1516), .Z(n_1517));
   INV_X1 i_839 (.A(n_1492), .ZN(n_1518));
   INV_X1 i_840 (.A(n_1473), .ZN(n_1519));
   AOI22_X1 i_841 (.A1(n_1518), .A2(n_1490), .B1(n_1519), .B2(n_1489), .ZN(
      n_1520));
   XNOR2_X1 i_842 (.A(n_1502), .B(n_1450), .ZN(n_1536));
   AOI22_X1 i_843 (.A1(n_1458), .A2(n_1463), .B1(n_1451), .B2(n_1457), .ZN(
      n_1537));
   OAI22_X1 i_844 (.A1(n_1433), .A2(n_1434), .B1(n_1375), .B2(n_1432), .ZN(
      n_1538));
   AOI21_X1 i_845 (.A(n_1319), .B1(n_1321), .B2(n_1323), .ZN(n_1539));
   XOR2_X1 i_846 (.A(n_1538), .B(n_1539), .Z(n_1540));
   OAI22_X1 i_847 (.A1(n_1437), .A2(n_1438), .B1(n_1344), .B2(n_1631), .ZN(
      n_1541));
   XNOR2_X1 i_848 (.A(n_1540), .B(n_1541), .ZN(n_1542));
   NAND2_X1 i_849 (.A1(n_1537), .A2(n_1542), .ZN(n_1543));
   OAI21_X1 i_850 (.A(n_1543), .B1(n_1537), .B2(n_1542), .ZN(n_1544));
   OAI22_X1 i_851 (.A1(n_1440), .A2(n_1445), .B1(n_1435), .B2(n_1439), .ZN(
      n_1545));
   XNOR2_X1 i_852 (.A(n_1544), .B(n_1545), .ZN(n_1546));
   XOR2_X1 i_853 (.A(n_1536), .B(n_1546), .Z(n_1547));
   INV_X1 i_854 (.A(n_1475), .ZN(n_1548));
   AOI22_X1 i_855 (.A1(n_1487), .A2(n_1488), .B1(n_1548), .B2(n_1486), .ZN(
      n_1549));
   XOR2_X1 i_856 (.A(n_1547), .B(n_1549), .Z(n_1550));
   INV_X1 i_857 (.A(n_1401), .ZN(n_1551));
   AOI22_X1 i_858 (.A1(n_1408), .A2(n_1416), .B1(n_1551), .B2(n_1407), .ZN(
      n_1552));
   XNOR2_X1 i_859 (.A(n_1616), .B(n_1615), .ZN(n_1556));
   OAI21_X1 i_860 (.A(n_1601), .B1(n_1604), .B2(n_1602), .ZN(n_1564));
   XOR2_X1 i_861 (.A(n_1556), .B(n_1564), .Z(n_1565));
   XOR2_X1 i_862 (.A(n_1587), .B(n_1508), .Z(n_1570));
   XOR2_X1 i_863 (.A(n_1565), .B(n_1570), .Z(n_1571));
   XNOR2_X1 i_864 (.A(n_1552), .B(n_1571), .ZN(n_1572));
   XOR2_X1 i_865 (.A(n_1636), .B(n_1635), .Z(n_1578));
   NAND3_X1 i_866 (.A1(n_1786), .A2(B[3]), .A3(A[21]), .ZN(n_1581));
   OAI22_X1 i_867 (.A1(n_1029), .A2(n_1317), .B1(n_424), .B2(n_1792), .ZN(n_1582));
   NAND2_X1 i_868 (.A1(n_1581), .A2(n_1582), .ZN(n_1583));
   XNOR2_X1 i_869 (.A(n_1583), .B(n_1318), .ZN(n_1584));
   XOR2_X1 i_870 (.A(n_1578), .B(n_1584), .Z(n_1585));
   XNOR2_X1 i_871 (.A(n_1627), .B(n_1626), .ZN(n_1591));
   XOR2_X1 i_872 (.A(n_1585), .B(n_1591), .Z(n_1592));
   XNOR2_X1 i_873 (.A(n_1572), .B(n_1592), .ZN(n_1593));
   XOR2_X1 i_874 (.A(n_1550), .B(n_1593), .Z(n_1594));
   XNOR2_X1 i_875 (.A(n_1520), .B(n_1594), .ZN(n_1595));
   XOR2_X1 i_876 (.A(n_1517), .B(n_1595), .Z(n_1596));
   XNOR2_X1 i_877 (.A(n_1500), .B(n_1596), .ZN(n_1597));
   XNOR2_X1 i_878 (.A(n_1498), .B(n_1597), .ZN(Out[26]));
   OAI22_X1 i_879 (.A1(n_1498), .A2(n_1597), .B1(n_1500), .B2(n_1596), .ZN(
      n_1598));
   INV_X1 i_880 (.A(n_1520), .ZN(n_1599));
   AOI22_X1 i_881 (.A1(n_1599), .A2(n_1594), .B1(n_1550), .B2(n_1593), .ZN(
      n_1600));
   XNOR2_X1 i_882 (.A(n_1655), .B(n_1658), .ZN(n_1618));
   OAI21_X1 i_883 (.A(n_1543), .B1(n_1544), .B2(n_1545), .ZN(n_1619));
   XNOR2_X1 i_884 (.A(n_1731), .B(n_1710), .ZN(n_1625));
   OAI21_X1 i_885 (.A(n_1745), .B1(n_1746), .B2(n_1791), .ZN(n_1632));
   XOR2_X1 i_886 (.A(n_1625), .B(n_1632), .Z(n_1633));
   XNOR2_X1 i_887 (.A(n_1612), .B(n_1611), .ZN(n_1637));
   XNOR2_X1 i_888 (.A(n_1633), .B(n_1637), .ZN(n_1638));
   XOR2_X1 i_889 (.A(n_1619), .B(n_1638), .Z(n_1639));
   XOR2_X1 i_890 (.A(n_1639), .B(n_1449), .Z(n_1641));
   XOR2_X1 i_891 (.A(n_1618), .B(n_1641), .Z(n_1642));
   INV_X1 i_892 (.A(n_1552), .ZN(n_1643));
   AOI22_X1 i_893 (.A1(n_1572), .A2(n_1592), .B1(n_1643), .B2(n_1571), .ZN(
      n_1644));
   XNOR2_X1 i_894 (.A(n_1642), .B(n_1644), .ZN(n_1645));
   XNOR2_X1 i_895 (.A(n_1600), .B(n_1645), .ZN(n_1646));
   XOR2_X1 i_896 (.A(n_1788), .B(n_1787), .Z(n_1651));
   XNOR2_X1 i_897 (.A(n_1762), .B(n_1648), .ZN(n_1656));
   XNOR2_X1 i_898 (.A(n_1651), .B(n_1656), .ZN(n_1657));
   XOR2_X1 i_899 (.A(n_1739), .B(n_1738), .Z(n_1663));
   OR2_X1 i_900 (.A1(n_1657), .A2(n_1663), .ZN(n_1664));
   INV_X1 i_901 (.A(n_1664), .ZN(n_1665));
   AOI21_X1 i_902 (.A(n_1665), .B1(n_1663), .B2(n_1657), .ZN(n_1666));
   XOR2_X1 i_903 (.A(n_1444), .B(n_1666), .Z(n_1667));
   AOI22_X1 i_904 (.A1(n_1509), .A2(n_1503), .B1(n_1521), .B2(n_1525), .ZN(
      n_1668));
   INV_X1 i_905 (.A(n_1541), .ZN(n_1669));
   INV_X1 i_906 (.A(n_1538), .ZN(n_1670));
   OAI22_X1 i_907 (.A1(n_1540), .A2(n_1669), .B1(n_1670), .B2(n_1539), .ZN(
      n_1671));
   XNOR2_X1 i_908 (.A(n_1668), .B(n_1671), .ZN(n_1672));
   OAI21_X1 i_909 (.A(n_1581), .B1(n_1583), .B2(n_1318), .ZN(n_1673));
   NOR2_X1 i_910 (.A1(n_340), .A2(n_1792), .ZN(n_1674));
   XOR2_X1 i_911 (.A(n_1673), .B(n_1674), .Z(n_1675));
   NOR2_X1 i_912 (.A1(n_1029), .A2(n_1881), .ZN(n_1677));
   XNOR2_X1 i_913 (.A(n_1675), .B(n_1677), .ZN(n_1678));
   XNOR2_X1 i_914 (.A(n_1672), .B(n_1678), .ZN(n_1679));
   AOI22_X1 i_915 (.A1(n_1565), .A2(n_1570), .B1(n_1556), .B2(n_1564), .ZN(
      n_1680));
   AOI22_X1 i_916 (.A1(n_1585), .A2(n_1591), .B1(n_1584), .B2(n_1578), .ZN(
      n_1681));
   XOR2_X1 i_917 (.A(n_1680), .B(n_1681), .Z(n_1682));
   XNOR2_X1 i_918 (.A(n_1679), .B(n_1682), .ZN(n_1683));
   XNOR2_X1 i_919 (.A(n_1667), .B(n_1683), .ZN(n_1684));
   INV_X1 i_920 (.A(n_1549), .ZN(n_1685));
   AOI22_X1 i_921 (.A1(n_1547), .A2(n_1685), .B1(n_1536), .B2(n_1546), .ZN(
      n_1686));
   XOR2_X1 i_922 (.A(n_1684), .B(n_1686), .Z(n_1687));
   INV_X1 i_923 (.A(n_1513), .ZN(n_1688));
   AOI22_X1 i_924 (.A1(n_1512), .A2(n_1688), .B1(n_1510), .B2(n_1511), .ZN(
      n_1689));
   XNOR2_X1 i_925 (.A(n_1687), .B(n_1689), .ZN(n_1690));
   XNOR2_X1 i_926 (.A(n_1646), .B(n_1690), .ZN(n_1691));
   AOI22_X1 i_927 (.A1(n_1517), .A2(n_1595), .B1(n_1516), .B2(n_1514), .ZN(
      n_1692));
   XOR2_X1 i_928 (.A(n_1691), .B(n_1692), .Z(n_1693));
   XNOR2_X1 i_929 (.A(n_1598), .B(n_1693), .ZN(Out[27]));
   AOI22_X1 i_930 (.A1(n_1598), .A2(n_1693), .B1(n_1691), .B2(n_1692), .ZN(
      n_1694));
   OAI22_X1 i_931 (.A1(n_1646), .A2(n_1690), .B1(n_1600), .B2(n_1645), .ZN(
      n_1695));
   XNOR2_X1 i_932 (.A(n_1694), .B(n_1695), .ZN(n_1696));
   AOI22_X1 i_933 (.A1(n_1687), .A2(n_1689), .B1(n_1684), .B2(n_1686), .ZN(
      n_1697));
   XNOR2_X1 i_934 (.A(n_1662), .B(n_1717), .ZN(n_1727));
   AOI22_X1 i_935 (.A1(n_1448), .A2(n_1639), .B1(n_1619), .B2(n_1638), .ZN(
      n_1729));
   XNOR2_X1 i_936 (.A(n_1734), .B(n_1730), .ZN(n_1735));
   XNOR2_X1 i_937 (.A(n_1825), .B(n_1573), .ZN(n_1741));
   XOR2_X1 i_938 (.A(n_1735), .B(n_1741), .Z(n_1742));
   XOR2_X1 i_939 (.A(n_1784), .B(n_1760), .Z(n_1747));
   XOR2_X1 i_940 (.A(n_1742), .B(n_1747), .Z(n_1748));
   XOR2_X1 i_941 (.A(n_1729), .B(n_1748), .Z(n_1749));
   XNOR2_X1 i_942 (.A(n_1727), .B(n_1749), .ZN(n_1750));
   XNOR2_X1 i_943 (.A(n_1697), .B(n_1750), .ZN(n_1751));
   AOI22_X1 i_944 (.A1(n_1679), .A2(n_1682), .B1(n_1681), .B2(n_1680), .ZN(
      n_1752));
   AOI22_X1 i_945 (.A1(n_1675), .A2(n_1677), .B1(n_1673), .B2(n_1674), .ZN(
      n_1753));
   NAND2_X1 i_946 (.A1(n_1893), .A2(n_1880), .ZN(n_1756));
   XNOR2_X1 i_947 (.A(n_1756), .B(n_1882), .ZN(n_1758));
   XNOR2_X1 i_948 (.A(n_1753), .B(n_1758), .ZN(n_1759));
   XOR2_X1 i_949 (.A(n_1877), .B(n_1878), .Z(n_1764));
   XNOR2_X1 i_950 (.A(n_1759), .B(n_1764), .ZN(n_1765));
   XOR2_X1 i_951 (.A(n_1752), .B(n_1765), .Z(n_1766));
   INV_X1 i_952 (.A(n_1671), .ZN(n_1767));
   AOI22_X1 i_953 (.A1(n_1672), .A2(n_1678), .B1(n_1668), .B2(n_1767), .ZN(
      n_1768));
   AOI22_X1 i_954 (.A1(n_1633), .A2(n_1637), .B1(n_1625), .B2(n_1632), .ZN(
      n_1769));
   OAI21_X1 i_955 (.A(n_1664), .B1(n_1656), .B2(n_1651), .ZN(n_1770));
   XNOR2_X1 i_956 (.A(n_1769), .B(n_1770), .ZN(n_1771));
   XNOR2_X1 i_957 (.A(n_1768), .B(n_1771), .ZN(n_1772));
   XNOR2_X1 i_958 (.A(n_1766), .B(n_1772), .ZN(n_1773));
   AOI22_X1 i_959 (.A1(n_1667), .A2(n_1683), .B1(n_1444), .B2(n_1666), .ZN(
      n_1774));
   XOR2_X1 i_960 (.A(n_1773), .B(n_1774), .Z(n_1775));
   INV_X1 i_961 (.A(n_1644), .ZN(n_1776));
   AOI22_X1 i_962 (.A1(n_1642), .A2(n_1776), .B1(n_1618), .B2(n_1641), .ZN(
      n_1777));
   XOR2_X1 i_963 (.A(n_1775), .B(n_1777), .Z(n_1778));
   XOR2_X1 i_964 (.A(n_1751), .B(n_1778), .Z(n_1779));
   XNOR2_X1 i_965 (.A(n_1696), .B(n_1779), .ZN(Out[28]));
   OAI22_X1 i_966 (.A1(n_1696), .A2(n_1779), .B1(n_1694), .B2(n_1695), .ZN(
      n_1780));
   AOI22_X1 i_967 (.A1(n_1775), .A2(n_1777), .B1(n_1773), .B2(n_1774), .ZN(
      n_1781));
   OAI21_X1 i_968 (.A(n_1891), .B1(n_1889), .B2(n_1890), .ZN(n_1798));
   XOR2_X1 i_969 (.A(n_1718), .B(n_1798), .Z(n_1799));
   INV_X1 i_970 (.A(n_1768), .ZN(n_1800));
   INV_X1 i_971 (.A(n_1769), .ZN(n_1801));
   AOI22_X1 i_972 (.A1(n_1800), .A2(n_1771), .B1(n_1801), .B2(n_1770), .ZN(
      n_1802));
   INV_X1 i_973 (.A(n_1753), .ZN(n_1803));
   AOI22_X1 i_974 (.A1(n_1759), .A2(n_1764), .B1(n_1803), .B2(n_1758), .ZN(
      n_1804));
   XOR2_X1 i_975 (.A(n_1804), .B(n_1719), .Z(n_1816));
   XNOR2_X1 i_976 (.A(n_1802), .B(n_1816), .ZN(n_1817));
   XNOR2_X1 i_977 (.A(n_1799), .B(n_1817), .ZN(n_1818));
   XNOR2_X1 i_978 (.A(n_1781), .B(n_1818), .ZN(n_1819));
   AOI22_X1 i_979 (.A1(n_1766), .A2(n_1772), .B1(n_1752), .B2(n_1765), .ZN(
      n_1820));
   AOI22_X1 i_980 (.A1(n_1742), .A2(n_1747), .B1(n_1735), .B2(n_1741), .ZN(
      n_1835));
   XNOR2_X1 i_981 (.A(n_1535), .B(n_1835), .ZN(n_1836));
   XOR2_X1 i_982 (.A(n_1806), .B(n_1805), .Z(n_1854));
   XNOR2_X1 i_983 (.A(n_1836), .B(n_1854), .ZN(n_1855));
   XOR2_X1 i_984 (.A(n_1820), .B(n_1855), .Z(n_1856));
   AOI22_X1 i_985 (.A1(n_1727), .A2(n_1749), .B1(n_1729), .B2(n_1748), .ZN(
      n_1857));
   XOR2_X1 i_986 (.A(n_1856), .B(n_1857), .Z(n_1858));
   XNOR2_X1 i_987 (.A(n_1819), .B(n_1858), .ZN(n_1859));
   INV_X1 i_988 (.A(n_1697), .ZN(n_1860));
   AOI22_X1 i_989 (.A1(n_1751), .A2(n_1778), .B1(n_1860), .B2(n_1750), .ZN(
      n_1861));
   XOR2_X1 i_990 (.A(n_1859), .B(n_1861), .Z(n_1862));
   XNOR2_X1 i_991 (.A(n_1780), .B(n_1862), .ZN(Out[29]));
   AOI22_X1 i_992 (.A1(n_1780), .A2(n_1862), .B1(n_1859), .B2(n_1861), .ZN(
      n_1863));
   INV_X1 i_993 (.A(n_1781), .ZN(n_1864));
   AOI22_X1 i_994 (.A1(n_1819), .A2(n_1858), .B1(n_1864), .B2(n_1818), .ZN(
      n_1865));
   INV_X1 i_995 (.A(n_1865), .ZN(n_1866));
   AOI22_X1 i_996 (.A1(n_1856), .A2(n_1857), .B1(n_1820), .B2(n_1855), .ZN(
      n_1867));
   INV_X1 i_997 (.A(n_1802), .ZN(n_1898));
   AOI22_X1 i_998 (.A1(n_1898), .A2(n_1816), .B1(n_1719), .B2(n_1804), .ZN(
      n_1899));
   XNOR2_X1 i_999 (.A(n_1793), .B(n_1899), .ZN(n_1900));
   XOR2_X1 i_1000 (.A(n_1867), .B(n_1900), .Z(n_1901));
   AOI22_X1 i_1001 (.A1(n_1799), .A2(n_1817), .B1(n_1718), .B2(n_1798), .ZN(
      n_1902));
   INV_X1 i_1002 (.A(n_1835), .ZN(n_1903));
   AOI22_X1 i_1003 (.A1(n_1836), .A2(n_1854), .B1(n_1535), .B2(n_1903), .ZN(
      n_1904));
   XNOR2_X1 i_1004 (.A(n_1935), .B(n_1931), .ZN(n_1919));
   XOR2_X1 i_1005 (.A(n_1914), .B(n_1910), .Z(n_1937));
   OR2_X1 i_1006 (.A1(n_1919), .A2(n_1937), .ZN(n_1938));
   NAND2_X1 i_1007 (.A1(n_1919), .A2(n_1937), .ZN(n_1939));
   NAND2_X1 i_1008 (.A1(n_1938), .A2(n_1939), .ZN(n_1940));
   XNOR2_X1 i_1009 (.A(n_1940), .B(n_1892), .ZN(n_1942));
   XNOR2_X1 i_1010 (.A(n_1904), .B(n_1942), .ZN(n_1943));
   XOR2_X1 i_1011 (.A(n_1902), .B(n_1943), .Z(n_1944));
   XNOR2_X1 i_1012 (.A(n_1901), .B(n_1944), .ZN(n_1945));
   NAND2_X1 i_1013 (.A1(n_1866), .A2(n_1945), .ZN(n_1946));
   OR2_X1 i_1014 (.A1(n_1945), .A2(n_1866), .ZN(n_1947));
   NAND2_X1 i_1015 (.A1(n_1946), .A2(n_1947), .ZN(n_1948));
   XNOR2_X1 i_1016 (.A(n_1863), .B(n_1948), .ZN(Out[30]));
   INV_X1 i_1017 (.A(n_1946), .ZN(n_1949));
   OAI21_X1 i_1018 (.A(n_1947), .B1(n_1863), .B2(n_1949), .ZN(n_1950));
   XOR2_X1 i_1019 (.A(n_2064), .B(n_2066), .Z(n_1968));
   INV_X1 i_1020 (.A(n_1938), .ZN(n_1969));
   AOI21_X1 i_1021 (.A(n_1969), .B1(n_1892), .B2(n_1939), .ZN(n_1970));
   XNOR2_X1 i_1022 (.A(n_1968), .B(n_1970), .ZN(n_1971));
   AOI22_X1 i_1023 (.A1(n_1793), .A2(n_1899), .B1(n_1812), .B2(n_1794), .ZN(
      n_1972));
   XOR2_X1 i_1024 (.A(n_1971), .B(n_1972), .Z(n_1973));
   XOR2_X1 i_1025 (.A(n_1895), .B(n_1930), .Z(n_1983));
   XNOR2_X1 i_1026 (.A(n_2119), .B(n_1964), .ZN(n_1989));
   XNOR2_X1 i_1027 (.A(n_2131), .B(n_2130), .ZN(n_1993));
   XOR2_X1 i_1028 (.A(n_1989), .B(n_1993), .Z(n_1994));
   NAND2_X1 i_1029 (.A1(A[13]), .A2(B[18]), .ZN(n_1995));
   XNOR2_X1 i_1030 (.A(n_1929), .B(n_1995), .ZN(n_1996));
   NAND2_X1 i_1031 (.A1(A[11]), .A2(B[20]), .ZN(n_1997));
   XNOR2_X1 i_1032 (.A(n_1996), .B(n_1997), .ZN(n_1998));
   XOR2_X1 i_1033 (.A(n_1994), .B(n_1998), .Z(n_1999));
   OR2_X1 i_1034 (.A1(n_1983), .A2(n_1999), .ZN(n_2000));
   NAND2_X1 i_1035 (.A1(n_1983), .A2(n_1999), .ZN(n_2001));
   NAND2_X1 i_1036 (.A1(n_2000), .A2(n_2001), .ZN(n_2002));
   XNOR2_X1 i_1037 (.A(n_1840), .B(n_2132), .ZN(n_2004));
   NAND2_X1 i_1038 (.A1(A[8]), .A2(B[23]), .ZN(n_2005));
   XNOR2_X1 i_1039 (.A(n_2004), .B(n_2005), .ZN(n_2006));
   INV_X1 i_1040 (.A(n_1821), .ZN(n_2007));
   AOI22_X1 i_1041 (.A1(n_1823), .A2(n_1814), .B1(n_2007), .B2(n_1815), .ZN(
      n_2008));
   XOR2_X1 i_1042 (.A(n_2006), .B(n_2008), .Z(n_2009));
   OAI33_X1 i_1043 (.A1(n_1912), .A2(n_558), .A3(n_560), .B1(n_1848), .B2(n_256), 
      .B3(n_1232), .ZN(n_2010));
   AOI21_X1 i_1044 (.A(n_1928), .B1(n_1926), .B2(n_1925), .ZN(n_2011));
   XNOR2_X1 i_1045 (.A(n_2010), .B(n_2011), .ZN(n_2012));
   AOI21_X1 i_1046 (.A(n_1837), .B1(n_1838), .B2(n_1841), .ZN(n_2013));
   XNOR2_X1 i_1047 (.A(n_2012), .B(n_2013), .ZN(n_2014));
   XNOR2_X1 i_1048 (.A(n_2009), .B(n_2014), .ZN(n_2015));
   XOR2_X1 i_1049 (.A(n_2002), .B(n_2015), .Z(n_2016));
   XOR2_X1 i_1050 (.A(n_1973), .B(n_2016), .Z(n_2017));
   OAI22_X1 i_1051 (.A1(n_1902), .A2(n_1943), .B1(n_1904), .B2(n_1942), .ZN(
      n_2018));
   XNOR2_X1 i_1052 (.A(n_2017), .B(n_2018), .ZN(n_2019));
   AOI22_X1 i_1053 (.A1(n_1901), .A2(n_1944), .B1(n_1867), .B2(n_1900), .ZN(
      n_2020));
   XOR2_X1 i_1054 (.A(n_2019), .B(n_2020), .Z(n_2021));
   NAND2_X1 i_1055 (.A1(n_1950), .A2(n_2021), .ZN(n_2022));
   OAI21_X1 i_1056 (.A(n_2022), .B1(n_1950), .B2(n_2021), .ZN(Out[31]));
   OAI21_X1 i_1057 (.A(n_2022), .B1(n_2020), .B2(n_2019), .ZN(n_2023));
   AOI22_X1 i_1058 (.A1(n_2017), .A2(n_2018), .B1(n_1973), .B2(n_2016), .ZN(
      n_2024));
   OAI21_X1 i_1059 (.A(n_2060), .B1(n_2053), .B2(n_2052), .ZN(n_2027));
   XOR2_X1 i_1060 (.A(n_1894), .B(n_2027), .Z(n_2028));
   AOI22_X1 i_1061 (.A1(n_2014), .A2(n_2009), .B1(n_2008), .B2(n_2006), .ZN(
      n_2029));
   XNOR2_X1 i_1062 (.A(n_2028), .B(n_2029), .ZN(n_2030));
   INV_X1 i_1063 (.A(n_2011), .ZN(n_2031));
   AOI22_X1 i_1064 (.A1(n_2012), .A2(n_2013), .B1(n_2010), .B2(n_2031), .ZN(
      n_2032));
   OAI22_X1 i_1065 (.A1(n_1996), .A2(n_1997), .B1(n_1929), .B2(n_1995), .ZN(
      n_2033));
   OAI22_X1 i_1066 (.A1(n_2004), .A2(n_2005), .B1(n_1840), .B2(n_2132), .ZN(
      n_2034));
   XNOR2_X1 i_1067 (.A(n_2033), .B(n_2034), .ZN(n_2035));
   XNOR2_X1 i_1068 (.A(n_2032), .B(n_2035), .ZN(n_2036));
   XNOR2_X1 i_1069 (.A(n_2125), .B(n_2118), .ZN(n_2042));
   XOR2_X1 i_1070 (.A(n_2036), .B(n_2042), .Z(n_2043));
   AOI22_X1 i_1071 (.A1(n_1994), .A2(n_1998), .B1(n_1989), .B2(n_1993), .ZN(
      n_2044));
   XNOR2_X1 i_1072 (.A(n_2043), .B(n_2044), .ZN(n_2045));
   INV_X1 i_1073 (.A(n_2000), .ZN(n_2046));
   OAI21_X1 i_1074 (.A(n_2001), .B1(n_2015), .B2(n_2046), .ZN(n_2047));
   OR2_X1 i_1075 (.A1(n_2045), .A2(n_2047), .ZN(n_2048));
   NAND2_X1 i_1076 (.A1(n_2045), .A2(n_2047), .ZN(n_2049));
   NAND2_X1 i_1077 (.A1(n_2048), .A2(n_2049), .ZN(n_2050));
   XNOR2_X1 i_1078 (.A(n_2030), .B(n_2050), .ZN(n_2051));
   XOR2_X1 i_1079 (.A(n_2068), .B(n_2071), .Z(n_2089));
   XOR2_X1 i_1080 (.A(n_2051), .B(n_2089), .Z(n_2090));
   INV_X1 i_1081 (.A(n_1972), .ZN(n_2091));
   INV_X1 i_1082 (.A(n_1970), .ZN(n_2092));
   AOI22_X1 i_1083 (.A1(n_1971), .A2(n_2091), .B1(n_1968), .B2(n_2092), .ZN(
      n_2093));
   XNOR2_X1 i_1084 (.A(n_2090), .B(n_2093), .ZN(n_2094));
   NOR2_X1 i_1085 (.A1(n_2024), .A2(n_2094), .ZN(n_2095));
   NAND2_X1 i_1086 (.A1(n_2024), .A2(n_2094), .ZN(n_2096));
   INV_X1 i_1087 (.A(n_2096), .ZN(n_2097));
   NOR2_X1 i_1088 (.A1(n_2095), .A2(n_2097), .ZN(n_2098));
   XNOR2_X1 i_1089 (.A(n_2023), .B(n_2098), .ZN(Out[32]));
   AOI21_X1 i_1090 (.A(n_2095), .B1(n_2023), .B2(n_2096), .ZN(n_2099));
   INV_X1 i_1091 (.A(n_2049), .ZN(n_2100));
   AOI21_X1 i_1092 (.A(n_2100), .B1(n_2030), .B2(n_2048), .ZN(n_2101));
   INV_X1 i_1093 (.A(n_2044), .ZN(n_2102));
   AOI22_X1 i_1094 (.A1(n_2043), .A2(n_2102), .B1(n_2036), .B2(n_2042), .ZN(
      n_2103));
   INV_X1 i_1095 (.A(n_2033), .ZN(n_2104));
   INV_X1 i_1096 (.A(n_2034), .ZN(n_2105));
   OAI22_X1 i_1097 (.A1(n_2032), .A2(n_2035), .B1(n_2104), .B2(n_2105), .ZN(
      n_2106));
   XOR2_X1 i_1098 (.A(n_2212), .B(n_2211), .Z(n_2112));
   XOR2_X1 i_1099 (.A(n_2106), .B(n_2112), .Z(n_2113));
   XOR2_X1 i_1100 (.A(n_2217), .B(n_2218), .Z(n_2120));
   XNOR2_X1 i_1101 (.A(n_2113), .B(n_2120), .ZN(n_2121));
   XOR2_X1 i_1102 (.A(n_2081), .B(n_2080), .Z(n_2138));
   XOR2_X1 i_1103 (.A(n_2121), .B(n_2138), .Z(n_2139));
   XOR2_X1 i_1104 (.A(n_2103), .B(n_2139), .Z(n_2140));
   XOR2_X1 i_1105 (.A(n_2101), .B(n_2140), .Z(n_2141));
   AOI22_X1 i_1106 (.A1(n_2028), .A2(n_2029), .B1(n_2027), .B2(n_1894), .ZN(
      n_2144));
   XOR2_X1 i_1107 (.A(n_2086), .B(n_2111), .Z(n_2155));
   AOI22_X1 i_1108 (.A1(n_1976), .A2(n_1981), .B1(n_1962), .B2(n_1975), .ZN(
      n_2156));
   XOR2_X1 i_1109 (.A(n_2155), .B(n_2156), .Z(n_2157));
   INV_X1 i_1110 (.A(n_1984), .ZN(n_2158));
   AOI22_X1 i_1111 (.A1(n_1991), .A2(n_2038), .B1(n_2158), .B2(n_1990), .ZN(
      n_2159));
   XOR2_X1 i_1112 (.A(n_2157), .B(n_2159), .Z(n_2160));
   XOR2_X1 i_1113 (.A(n_2144), .B(n_2160), .Z(n_2161));
   XNOR2_X1 i_1114 (.A(n_2073), .B(n_2161), .ZN(n_2162));
   XOR2_X1 i_1115 (.A(n_2141), .B(n_2162), .Z(n_2163));
   AOI22_X1 i_1116 (.A1(n_2093), .A2(n_2090), .B1(n_2089), .B2(n_2051), .ZN(
      n_2164));
   OR2_X1 i_1117 (.A1(n_2163), .A2(n_2164), .ZN(n_2165));
   NAND2_X1 i_1118 (.A1(n_2163), .A2(n_2164), .ZN(n_2166));
   NAND2_X1 i_1119 (.A1(n_2165), .A2(n_2166), .ZN(n_2167));
   XNOR2_X1 i_1120 (.A(n_2099), .B(n_2167), .ZN(Out[33]));
   INV_X1 i_1121 (.A(n_2166), .ZN(n_2168));
   AOI21_X1 i_1122 (.A(n_2168), .B1(n_2099), .B2(n_2165), .ZN(n_2169));
   AOI22_X1 i_1123 (.A1(n_2141), .A2(n_2162), .B1(n_2140), .B2(n_2101), .ZN(
      n_2170));
   AOI22_X1 i_1124 (.A1(n_2073), .A2(n_2161), .B1(n_2144), .B2(n_2160), .ZN(
      n_2171));
   XNOR2_X1 i_1125 (.A(n_2194), .B(n_2179), .ZN(n_2189));
   AOI22_X1 i_1126 (.A1(n_2113), .A2(n_2120), .B1(n_2106), .B2(n_2112), .ZN(
      n_2190));
   XOR2_X1 i_1127 (.A(n_2189), .B(n_2190), .Z(n_2191));
   INV_X1 i_1128 (.A(n_2110), .ZN(n_2192));
   AOI22_X1 i_1129 (.A1(n_2107), .A2(n_2087), .B1(n_2192), .B2(n_2109), .ZN(
      n_2193));
   XOR2_X1 i_1130 (.A(n_2246), .B(n_2248), .Z(n_2197));
   XNOR2_X1 i_1131 (.A(n_2193), .B(n_2197), .ZN(n_2198));
   XOR2_X1 i_1132 (.A(n_2253), .B(n_2256), .Z(n_2203));
   XNOR2_X1 i_1133 (.A(n_2198), .B(n_2203), .ZN(n_2204));
   XOR2_X1 i_1134 (.A(n_2191), .B(n_2204), .Z(n_2205));
   XNOR2_X1 i_1135 (.A(n_2171), .B(n_2205), .ZN(n_2206));
   INV_X1 i_1136 (.A(n_2103), .ZN(n_2207));
   AOI22_X1 i_1137 (.A1(n_2139), .A2(n_2207), .B1(n_2121), .B2(n_2138), .ZN(
      n_2208));
   XOR2_X1 i_1138 (.A(n_2085), .B(n_2076), .Z(n_2219));
   INV_X1 i_1139 (.A(n_2159), .ZN(n_2220));
   AOI22_X1 i_1140 (.A1(n_2157), .A2(n_2220), .B1(n_2155), .B2(n_2156), .ZN(
      n_2221));
   XOR2_X1 i_1141 (.A(n_2219), .B(n_2221), .Z(n_2222));
   XNOR2_X1 i_1142 (.A(n_2208), .B(n_2222), .ZN(n_2223));
   XOR2_X1 i_1143 (.A(n_2206), .B(n_2223), .Z(n_2224));
   XOR2_X1 i_1144 (.A(n_2170), .B(n_2224), .Z(n_2225));
   XNOR2_X1 i_1145 (.A(n_2169), .B(n_2225), .ZN(Out[34]));
   AOI22_X1 i_1146 (.A1(n_2169), .A2(n_2225), .B1(n_2224), .B2(n_2170), .ZN(
      n_2226));
   INV_X1 i_1147 (.A(n_2208), .ZN(n_2227));
   AOI22_X1 i_1148 (.A1(n_2227), .A2(n_2222), .B1(n_2221), .B2(n_2219), .ZN(
      n_2228));
   AOI22_X1 i_1149 (.A1(n_2191), .A2(n_2204), .B1(n_2190), .B2(n_2189), .ZN(
      n_2229));
   INV_X1 i_1150 (.A(n_2216), .ZN(n_2230));
   INV_X1 i_1151 (.A(n_2196), .ZN(n_2231));
   AOI22_X1 i_1152 (.A1(n_2230), .A2(n_2195), .B1(n_2210), .B2(n_2231), .ZN(
      n_2232));
   XNOR2_X1 i_1153 (.A(n_2260), .B(n_2261), .ZN(n_2237));
   XOR2_X1 i_1154 (.A(n_2232), .B(n_2237), .Z(n_2238));
   INV_X1 i_1155 (.A(n_2193), .ZN(n_2239));
   AOI22_X1 i_1156 (.A1(n_2198), .A2(n_2203), .B1(n_2239), .B2(n_2197), .ZN(
      n_2240));
   XNOR2_X1 i_1157 (.A(n_2238), .B(n_2240), .ZN(n_2241));
   XNOR2_X1 i_1158 (.A(n_2496), .B(n_2495), .ZN(n_2247));
   XNOR2_X1 i_1159 (.A(n_2501), .B(n_2500), .ZN(n_2254));
   XOR2_X1 i_1160 (.A(n_2247), .B(n_2254), .Z(n_2255));
   XNOR2_X1 i_1161 (.A(n_2486), .B(n_2485), .ZN(n_2262));
   XNOR2_X1 i_1162 (.A(n_2255), .B(n_2262), .ZN(n_2263));
   XOR2_X1 i_1163 (.A(n_2241), .B(n_2263), .Z(n_2264));
   XNOR2_X1 i_1164 (.A(n_2229), .B(n_2264), .ZN(n_2265));
   XOR2_X1 i_1165 (.A(n_2265), .B(n_2074), .Z(n_2282));
   XOR2_X1 i_1166 (.A(n_2228), .B(n_2282), .Z(n_2283));
   INV_X1 i_1167 (.A(n_2171), .ZN(n_2284));
   AOI22_X1 i_1168 (.A1(n_2206), .A2(n_2223), .B1(n_2284), .B2(n_2205), .ZN(
      n_2285));
   OR2_X1 i_1169 (.A1(n_2283), .A2(n_2285), .ZN(n_2286));
   NAND2_X1 i_1170 (.A1(n_2283), .A2(n_2285), .ZN(n_2287));
   NAND2_X1 i_1171 (.A1(n_2286), .A2(n_2287), .ZN(n_2288));
   XNOR2_X1 i_1172 (.A(n_2226), .B(n_2288), .ZN(Out[35]));
   INV_X1 i_1173 (.A(n_2287), .ZN(n_2289));
   AOI21_X1 i_1174 (.A(n_2289), .B1(n_2226), .B2(n_2286), .ZN(n_2290));
   INV_X1 i_1175 (.A(n_2228), .ZN(n_2291));
   AOI22_X1 i_1176 (.A1(n_2282), .A2(n_2291), .B1(n_2265), .B2(n_2074), .ZN(
      n_2292));
   AOI22_X1 i_1177 (.A1(n_2229), .A2(n_2264), .B1(n_2241), .B2(n_2263), .ZN(
      n_2293));
   AOI22_X1 i_1178 (.A1(n_2238), .A2(n_2240), .B1(n_2232), .B2(n_2237), .ZN(
      n_2294));
   AOI22_X1 i_1179 (.A1(n_2146), .A2(n_2135), .B1(n_2148), .B2(n_2147), .ZN(
      n_2295));
   AOI22_X1 i_1180 (.A1(n_2255), .A2(n_2262), .B1(n_2247), .B2(n_2254), .ZN(
      n_2296));
   XNOR2_X1 i_1181 (.A(n_2295), .B(n_2296), .ZN(n_2297));
   XOR2_X1 i_1182 (.A(n_2294), .B(n_2297), .Z(n_2298));
   XNOR2_X1 i_1183 (.A(n_2293), .B(n_2298), .ZN(n_2299));
   INV_X1 i_1184 (.A(n_2178), .ZN(n_2300));
   AOI22_X1 i_1185 (.A1(n_2133), .A2(n_2075), .B1(n_2300), .B2(n_2134), .ZN(
      n_2301));
   INV_X1 i_1186 (.A(n_2275), .ZN(n_2313));
   NAND2_X1 i_1187 (.A1(n_2313), .A2(n_2281), .ZN(n_2315));
   XNOR2_X1 i_1188 (.A(n_2315), .B(n_2280), .ZN(n_2321));
   XNOR2_X1 i_1189 (.A(n_2490), .B(n_2484), .ZN(n_2328));
   XNOR2_X1 i_1190 (.A(n_2481), .B(n_2480), .ZN(n_2334));
   OAI21_X1 i_1191 (.A(n_2457), .B1(n_2458), .B2(n_2506), .ZN(n_2342));
   XOR2_X1 i_1192 (.A(n_2334), .B(n_2342), .Z(n_2343));
   NAND2_X1 i_1193 (.A1(n_2328), .A2(n_2343), .ZN(n_2344));
   OAI21_X1 i_1194 (.A(n_2344), .B1(n_2343), .B2(n_2328), .ZN(n_2345));
   XOR2_X1 i_1195 (.A(n_2321), .B(n_2345), .Z(n_2346));
   XNOR2_X1 i_1196 (.A(n_2301), .B(n_2346), .ZN(n_2347));
   XNOR2_X1 i_1197 (.A(n_2299), .B(n_2347), .ZN(n_2348));
   XNOR2_X1 i_1198 (.A(n_2292), .B(n_2348), .ZN(n_2349));
   XNOR2_X1 i_2386 (.A(n_2290), .B(n_2349), .ZN(Out[36]));
   INV_X1 i_1199 (.A(n_2292), .ZN(n_2350));
   AOI22_X1 i_1200 (.A1(n_2290), .A2(n_2349), .B1(n_2350), .B2(n_2348), .ZN(
      n_2351));
   AOI22_X1 i_1201 (.A1(n_2301), .A2(n_2346), .B1(n_2321), .B2(n_2345), .ZN(
      n_2352));
   XNOR2_X1 i_1202 (.A(n_2455), .B(n_2454), .ZN(n_2358));
   XNOR2_X1 i_1203 (.A(n_2302), .B(n_2358), .ZN(n_2359));
   XNOR2_X1 i_1204 (.A(n_2467), .B(n_2466), .ZN(n_2365));
   XOR2_X1 i_1205 (.A(n_2359), .B(n_2365), .Z(n_2366));
   XOR2_X1 i_1206 (.A(n_2352), .B(n_2366), .Z(n_2367));
   INV_X1 i_1207 (.A(n_2295), .ZN(n_2368));
   AOI22_X1 i_1208 (.A1(n_2294), .A2(n_2297), .B1(n_2368), .B2(n_2296), .ZN(
      n_2369));
   XOR2_X1 i_1209 (.A(n_2336), .B(n_2335), .Z(n_2375));
   XOR2_X1 i_1210 (.A(n_2326), .B(n_2325), .Z(n_2379));
   XOR2_X1 i_1211 (.A(n_2375), .B(n_2379), .Z(n_2380));
   XOR2_X1 i_1212 (.A(n_2341), .B(n_2340), .Z(n_2385));
   XNOR2_X1 i_1213 (.A(n_2380), .B(n_2385), .ZN(n_2386));
   OAI21_X1 i_1214 (.A(n_2344), .B1(n_2342), .B2(n_2334), .ZN(n_2387));
   XOR2_X1 i_1215 (.A(n_2386), .B(n_2387), .Z(n_2388));
   XNOR2_X1 i_1216 (.A(n_2369), .B(n_2388), .ZN(n_2389));
   XOR2_X1 i_1217 (.A(n_2367), .B(n_2389), .Z(n_2390));
   INV_X1 i_1218 (.A(n_2293), .ZN(n_2391));
   AOI22_X1 i_1219 (.A1(n_2299), .A2(n_2347), .B1(n_2391), .B2(n_2298), .ZN(
      n_2392));
   XOR2_X1 i_1220 (.A(n_2390), .B(n_2392), .Z(n_2393));
   XNOR2_X1 i_2431 (.A(n_2351), .B(n_2393), .ZN(Out[37]));
   INV_X1 i_1221 (.A(n_2392), .ZN(n_2394));
   OAI22_X1 i_1222 (.A1(n_2351), .A2(n_2393), .B1(n_2394), .B2(n_2390), .ZN(
      n_2395));
   INV_X1 i_1223 (.A(n_2352), .ZN(n_2396));
   OAI22_X1 i_1224 (.A1(n_2367), .A2(n_2389), .B1(n_2396), .B2(n_2366), .ZN(
      n_2397));
   INV_X1 i_1225 (.A(n_2387), .ZN(n_2398));
   OAI22_X1 i_1226 (.A1(n_2369), .A2(n_2388), .B1(n_2398), .B2(n_2386), .ZN(
      n_2399));
   AOI22_X1 i_1227 (.A1(n_2359), .A2(n_2365), .B1(n_2303), .B2(n_2358), .ZN(
      n_2401));
   XOR2_X1 i_1228 (.A(n_2399), .B(n_2401), .Z(n_2402));
   XOR2_X1 i_1229 (.A(n_2450), .B(n_2449), .Z(n_2414));
   AOI22_X1 i_1230 (.A1(n_2380), .A2(n_2385), .B1(n_2375), .B2(n_2379), .ZN(
      n_2415));
   XOR2_X1 i_1231 (.A(n_2414), .B(n_2415), .Z(n_2416));
   XNOR2_X1 i_1232 (.A(n_2462), .B(n_2461), .ZN(n_2434));
   XNOR2_X1 i_1233 (.A(n_2416), .B(n_2434), .ZN(n_2435));
   XOR2_X1 i_1234 (.A(n_2402), .B(n_2435), .Z(n_2436));
   NOR2_X1 i_1235 (.A1(n_2397), .A2(n_2436), .ZN(n_2437));
   NAND2_X1 i_1236 (.A1(n_2397), .A2(n_2436), .ZN(n_2438));
   INV_X1 i_2477 (.A(n_2438), .ZN(n_2439));
   NOR2_X1 i_2478 (.A1(n_2437), .A2(n_2439), .ZN(n_2440));
   XNOR2_X1 i_2479 (.A(n_2395), .B(n_2440), .ZN(Out[38]));
   AOI21_X1 i_1237 (.A(n_2437), .B1(n_2395), .B2(n_2438), .ZN(n_2441));
   XNOR2_X1 i_1238 (.A(n_2460), .B(n_2445), .ZN(n_2452));
   XOR2_X1 i_1239 (.A(n_2417), .B(n_2407), .Z(n_2470));
   XOR2_X1 i_1240 (.A(n_2452), .B(n_2470), .Z(n_2471));
   AOI22_X1 i_1241 (.A1(n_2434), .A2(n_2416), .B1(n_2414), .B2(n_2415), .ZN(
      n_2472));
   XNOR2_X1 i_1242 (.A(n_2471), .B(n_2472), .ZN(n_2473));
   XNOR2_X1 i_1243 (.A(n_2441), .B(n_2473), .ZN(n_2474));
   AOI22_X1 i_1244 (.A1(n_2402), .A2(n_2435), .B1(n_2399), .B2(n_2401), .ZN(
      n_2475));
   XNOR2_X1 i_2515 (.A(n_2474), .B(n_2475), .ZN(Out[39]));
   INV_X1 i_1245 (.A(n_2441), .ZN(n_2476));
   AOI22_X1 i_1246 (.A1(n_2474), .A2(n_2475), .B1(n_2476), .B2(n_2473), .ZN(
      n_2477));
   AOI22_X1 i_1247 (.A1(n_2471), .A2(n_2472), .B1(n_2452), .B2(n_2470), .ZN(
      n_2478));
   XNOR2_X1 i_1248 (.A(n_2444), .B(n_2382), .ZN(n_2509));
   XOR2_X1 i_1249 (.A(n_2478), .B(n_2509), .Z(n_2510));
   XOR2_X1 i_2551 (.A(n_2477), .B(n_2510), .Z(Out[40]));
   INV_X1 i_1250 (.A(n_2477), .ZN(n_2511));
   AOI22_X1 i_1251 (.A1(n_2511), .A2(n_2510), .B1(n_2478), .B2(n_2509), .ZN(
      n_2512));
   AOI22_X1 i_1252 (.A1(n_2444), .A2(n_2382), .B1(n_2405), .B2(n_2383), .ZN(
      n_2513));
   INV_X1 i_1253 (.A(n_2423), .ZN(n_2514));
   AOI21_X1 i_1254 (.A(n_2428), .B1(n_2514), .B2(n_2427), .ZN(n_2515));
   XOR2_X1 i_1255 (.A(n_2515), .B(n_2357), .Z(n_2522));
   XOR2_X1 i_1256 (.A(n_2587), .B(n_2370), .Z(n_2527));
   OAI21_X1 i_1257 (.A(n_2528), .B1(n_2526), .B2(n_2521), .ZN(n_2534));
   NOR2_X1 i_1258 (.A1(n_2527), .A2(n_2534), .ZN(n_2535));
   AOI21_X1 i_1259 (.A(n_2535), .B1(n_2534), .B2(n_2527), .ZN(n_2536));
   XNOR2_X1 i_1260 (.A(n_2522), .B(n_2536), .ZN(n_2537));
   AOI22_X1 i_1261 (.A1(n_2400), .A2(n_2384), .B1(n_2403), .B2(n_2404), .ZN(
      n_2538));
   XOR2_X1 i_1262 (.A(n_2537), .B(n_2538), .Z(n_2539));
   INV_X1 i_1263 (.A(n_2406), .ZN(n_2540));
   AOI22_X1 i_1264 (.A1(n_2420), .A2(n_2540), .B1(n_2421), .B2(n_2304), .ZN(
      n_2542));
   XOR2_X1 i_1265 (.A(n_2539), .B(n_2542), .Z(n_2543));
   NOR2_X1 i_1266 (.A1(n_2513), .A2(n_2543), .ZN(n_2544));
   NAND2_X1 i_1267 (.A1(n_2513), .A2(n_2543), .ZN(n_2545));
   INV_X1 i_2587 (.A(n_2545), .ZN(n_2546));
   NOR2_X1 i_2588 (.A1(n_2544), .A2(n_2546), .ZN(n_2547));
   XOR2_X1 i_2589 (.A(n_2512), .B(n_2547), .Z(Out[41]));
   AOI21_X1 i_1268 (.A(n_2544), .B1(n_2512), .B2(n_2545), .ZN(n_2548));
   AOI22_X1 i_2591 (.A1(n_2539), .A2(n_2542), .B1(n_2537), .B2(n_2538), .ZN(
      n_2549));
   INV_X1 i_2592 (.A(n_2549), .ZN(n_2550));
   OR2_X1 i_2593 (.A1(n_2548), .A2(n_2550), .ZN(n_2551));
   NAND2_X1 i_2594 (.A1(n_2548), .A2(n_2550), .ZN(n_2552));
   NAND2_X1 i_2595 (.A1(n_2551), .A2(n_2552), .ZN(n_2553));
   XNOR2_X1 i_2614 (.A(n_2590), .B(n_2584), .ZN(n_2572));
   AOI22_X1 i_2615 (.A1(n_2515), .A2(n_2357), .B1(n_2371), .B2(n_2360), .ZN(
      n_2573));
   XOR2_X1 i_2616 (.A(n_2572), .B(n_2573), .Z(n_2574));
   AOI21_X1 i_2617 (.A(n_2535), .B1(n_2522), .B2(n_2536), .ZN(n_2575));
   XNOR2_X1 i_2618 (.A(n_2574), .B(n_2575), .ZN(n_2576));
   XNOR2_X1 i_2619 (.A(n_2553), .B(n_2576), .ZN(Out[42]));
   INV_X1 i_2620 (.A(n_2551), .ZN(n_2577));
   OAI21_X1 i_2621 (.A(n_2552), .B1(n_2577), .B2(n_2576), .ZN(n_2578));
   AOI22_X1 i_2622 (.A1(n_2574), .A2(n_2575), .B1(n_2572), .B2(n_2573), .ZN(
      n_2579));
   XNOR2_X1 i_2637 (.A(n_2592), .B(n_2583), .ZN(n_2594));
   XNOR2_X1 i_2638 (.A(n_2579), .B(n_2594), .ZN(n_2595));
   XNOR2_X1 i_2639 (.A(n_2578), .B(n_2595), .ZN(Out[43]));
   INV_X1 i_2640 (.A(n_2579), .ZN(n_2596));
   AOI22_X1 i_2641 (.A1(n_2578), .A2(n_2595), .B1(n_2594), .B2(n_2596), .ZN(
      n_2597));
   INV_X1 i_2653 (.A(n_2580), .ZN(n_0));
   NOR2_X1 i_2654 (.A1(n_2582), .A2(n_2581), .ZN(n_1));
   NOR2_X1 i_2655 (.A1(n_0), .A2(n_1), .ZN(n_2));
   XOR2_X1 i_2656 (.A(n_2597), .B(n_2), .Z(Out[44]));
   INV_X1 i_2657 (.A(n_2597), .ZN(n_4));
   AOI21_X1 i_2658 (.A(n_1), .B1(n_4), .B2(n_2580), .ZN(n_5));
   OAI22_X1 i_1269 (.A1(n_2520), .A2(n_2562), .B1(n_2517), .B2(n_2519), .ZN(n_6));
   NAND2_X1 i_1270 (.A1(B[23]), .A2(A[23]), .ZN(n_7));
   NOR2_X1 i_1271 (.A1(n_2517), .A2(n_7), .ZN(n_8));
   AOI22_X1 i_1272 (.A1(A[22]), .A2(B[23]), .B1(B[22]), .B2(A[23]), .ZN(n_9));
   NOR2_X1 i_1273 (.A1(n_8), .A2(n_9), .ZN(n_10));
   XNOR2_X1 i_1274 (.A(n_6), .B(n_10), .ZN(n_11));
   XOR2_X1 i_2666 (.A(n_2569), .B(n_11), .Z(n_12));
   XNOR2_X1 i_2667 (.A(n_5), .B(n_12), .ZN(Out[45]));
   AOI21_X1 i_1275 (.A(n_11), .B1(n_2580), .B2(n_2570), .ZN(n_13));
   AOI21_X1 i_2670 (.A(n_1), .B1(n_2570), .B2(n_11), .ZN(n_14));
   AOI21_X1 i_2671 (.A(n_13), .B1(n_2597), .B2(n_14), .ZN(n_15));
   AOI21_X1 i_2672 (.A(n_8), .B1(n_6), .B2(n_10), .ZN(n_16));
   XOR2_X1 i_2673 (.A(n_16), .B(n_7), .Z(n_17));
   XNOR2_X1 i_2674 (.A(n_15), .B(n_17), .ZN(Out[46]));
   AOI21_X1 i_2675 (.A(n_7), .B1(n_15), .B2(n_17), .ZN(Out[47]));
   XNOR2_X1 i_1276 (.A(n_19), .B(n_18), .ZN(Out[2]));
   NAND2_X1 i_1277 (.A1(n_22), .A2(n_21), .ZN(n_18));
   NOR2_X1 i_1278 (.A1(n_27), .A2(n_20), .ZN(n_19));
   NAND2_X1 i_1279 (.A1(A[0]), .A2(B[0]), .ZN(n_20));
   OR2_X1 i_1280 (.A1(n_24), .A2(n_23), .ZN(n_21));
   NAND2_X1 i_1281 (.A1(n_24), .A2(n_23), .ZN(n_22));
   NOR2_X1 i_1282 (.A1(n_33), .A2(n_28), .ZN(n_23));
   AOI21_X1 i_1283 (.A(n_25), .B1(n_27), .B2(n_26), .ZN(n_24));
   NOR2_X1 i_1284 (.A1(n_27), .A2(n_26), .ZN(n_25));
   NAND2_X1 i_1285 (.A1(A[0]), .A2(B[2]), .ZN(n_26));
   NAND2_X1 i_1286 (.A1(A[1]), .A2(B[1]), .ZN(n_27));
   INV_X1 i_1287 (.A(B[0]), .ZN(n_28));
   INV_X1 i_1288 (.A(B[2]), .ZN(n_29));
   INV_X1 i_1289 (.A(A[0]), .ZN(n_31));
   INV_X1 i_1290 (.A(A[2]), .ZN(n_33));
   NAND2_X1 i_1291 (.A1(A[0]), .A2(B[3]), .ZN(n_64));
   AOI22_X1 i_1292 (.A1(A[1]), .A2(B[2]), .B1(A[2]), .B2(B[1]), .ZN(n_66));
   INV_X1 i_1293 (.A(A[3]), .ZN(n_99));
   NOR2_X1 i_1294 (.A1(n_99), .A2(n_28), .ZN(n_107));
   XNOR2_X1 i_1295 (.A(n_107), .B(n_25), .ZN(n_113));
   INV_X1 i_1296 (.A(n_22), .ZN(n_139));
   AOI21_X1 i_1297 (.A(n_139), .B1(n_19), .B2(n_21), .ZN(n_140));
   NOR2_X1 i_1298 (.A1(n_113), .A2(n_140), .ZN(n_141));
   INV_X1 i_1299 (.A(n_141), .ZN(n_142));
   NAND2_X1 i_1300 (.A1(n_113), .A2(n_140), .ZN(n_143));
   NAND2_X1 i_1301 (.A1(n_142), .A2(n_143), .ZN(n_146));
   NOR3_X1 i_1302 (.A1(n_27), .A2(n_33), .A3(n_29), .ZN(n_147));
   NOR2_X1 i_1303 (.A1(n_66), .A2(n_147), .ZN(n_148));
   XNOR2_X1 i_1304 (.A(n_148), .B(n_64), .ZN(n_149));
   XNOR2_X1 i_1305 (.A(n_146), .B(n_149), .ZN(Out[3]));
   INV_X1 i_1306 (.A(n_147), .ZN(n_150));
   NAND2_X1 i_1307 (.A1(B[5]), .A2(A[7]), .ZN(n_151));
   NAND2_X1 i_1308 (.A1(A[8]), .A2(B[4]), .ZN(n_166));
   NOR2_X1 i_1309 (.A1(n_151), .A2(n_166), .ZN(n_167));
   AOI21_X1 i_1310 (.A(n_167), .B1(n_151), .B2(n_166), .ZN(n_168));
   INV_X1 i_1311 (.A(B[6]), .ZN(n_169));
   INV_X1 i_1312 (.A(A[6]), .ZN(n_170));
   NOR2_X1 i_1313 (.A1(n_169), .A2(n_170), .ZN(n_171));
   NAND2_X1 i_1314 (.A1(n_168), .A2(n_171), .ZN(n_174));
   NAND2_X1 i_1315 (.A1(B[7]), .A2(A[5]), .ZN(n_175));
   NAND2_X1 i_1316 (.A1(B[8]), .A2(A[4]), .ZN(n_176));
   XNOR2_X1 i_1317 (.A(n_175), .B(n_176), .ZN(n_177));
   NAND2_X1 i_1318 (.A1(B[9]), .A2(A[3]), .ZN(n_178));
   INV_X1 i_1319 (.A(n_167), .ZN(n_181));
   NAND2_X1 i_1320 (.A1(n_174), .A2(n_181), .ZN(n_182));
   OAI22_X1 i_1321 (.A1(n_177), .A2(n_178), .B1(n_175), .B2(n_176), .ZN(n_187));
   NAND2_X1 i_1322 (.A1(n_182), .A2(n_187), .ZN(n_188));
   OAI21_X1 i_1323 (.A(n_188), .B1(n_182), .B2(n_187), .ZN(n_189));
   NAND2_X1 i_1324 (.A1(A[0]), .A2(B[11]), .ZN(n_198));
   NAND2_X1 i_1325 (.A1(B[12]), .A2(A[1]), .ZN(n_204));
   NOR2_X1 i_1326 (.A1(n_198), .A2(n_204), .ZN(n_205));
   AOI22_X1 i_1327 (.A1(B[12]), .A2(A[0]), .B1(A[1]), .B2(B[11]), .ZN(n_206));
   NOR2_X1 i_1328 (.A1(n_205), .A2(n_206), .ZN(n_207));
   NAND2_X1 i_1329 (.A1(B[10]), .A2(A[2]), .ZN(n_208));
   INV_X1 i_1330 (.A(n_208), .ZN(n_209));
   AOI21_X1 i_1331 (.A(n_205), .B1(n_207), .B2(n_209), .ZN(n_212));
   OAI21_X1 i_1332 (.A(n_188), .B1(n_189), .B2(n_212), .ZN(n_222));
   NAND2_X1 i_1333 (.A1(B[11]), .A2(A[2]), .ZN(n_226));
   NOR2_X1 i_1334 (.A1(n_204), .A2(n_226), .ZN(n_227));
   AOI21_X1 i_1335 (.A(n_227), .B1(n_204), .B2(n_226), .ZN(n_228));
   INV_X1 i_1336 (.A(B[13]), .ZN(n_229));
   NOR2_X1 i_1337 (.A1(n_229), .A2(n_31), .ZN(n_230));
   AOI21_X1 i_1338 (.A(n_227), .B1(n_228), .B2(n_230), .ZN(n_245));
   XNOR2_X1 i_1339 (.A(n_222), .B(n_245), .ZN(n_246));
   INV_X1 i_1340 (.A(A[13]), .ZN(n_256));
   INV_X1 i_1341 (.A(B[1]), .ZN(n_257));
   INV_X1 i_1342 (.A(A[12]), .ZN(n_258));
   OAI22_X1 i_1343 (.A1(n_258), .A2(n_257), .B1(n_256), .B2(n_28), .ZN(n_259));
   NAND2_X1 i_1344 (.A1(B[1]), .A2(A[11]), .ZN(n_260));
   NAND2_X1 i_1345 (.A1(B[2]), .A2(A[10]), .ZN(n_261));
   XNOR2_X1 i_1346 (.A(n_260), .B(n_261), .ZN(n_262));
   NAND2_X1 i_1347 (.A1(B[3]), .A2(A[9]), .ZN(n_263));
   OAI22_X1 i_1348 (.A1(n_262), .A2(n_263), .B1(n_260), .B2(n_261), .ZN(n_264));
   OR4_X1 i_1349 (.A1(n_256), .A2(n_258), .A3(n_257), .A4(n_28), .ZN(n_265));
   INV_X1 i_1350 (.A(n_265), .ZN(n_266));
   OAI21_X1 i_1351 (.A(n_259), .B1(n_264), .B2(n_266), .ZN(n_267));
   XNOR2_X1 i_1352 (.A(n_246), .B(n_267), .ZN(n_268));
   NOR2_X1 i_1353 (.A1(n_258), .A2(n_28), .ZN(n_269));
   NAND2_X1 i_1354 (.A1(B[5]), .A2(A[8]), .ZN(n_270));
   NAND2_X1 i_1355 (.A1(B[4]), .A2(A[7]), .ZN(n_272));
   XNOR2_X1 i_1356 (.A(n_304), .B(n_274), .ZN(n_273));
   AOI22_X1 i_1357 (.A1(n_279), .A2(n_277), .B1(n_276), .B2(n_275), .ZN(n_274));
   XNOR2_X1 i_1358 (.A(n_228), .B(n_230), .ZN(n_275));
   XOR2_X1 i_1359 (.A(n_279), .B(n_277), .Z(n_276));
   XOR2_X1 i_1360 (.A(n_270), .B(n_278), .Z(n_277));
   NOR2_X1 i_1361 (.A1(n_282), .A2(n_281), .ZN(n_278));
   XOR2_X1 i_1362 (.A(n_284), .B(n_280), .Z(n_279));
   NOR2_X1 i_1363 (.A1(n_286), .A2(n_285), .ZN(n_280));
   AOI22_X1 i_1364 (.A1(B[6]), .A2(A[7]), .B1(B[7]), .B2(A[6]), .ZN(n_281));
   INV_X1 i_1365 (.A(n_283), .ZN(n_282));
   NAND3_X1 i_1366 (.A1(A[7]), .A2(n_171), .A3(B[7]), .ZN(n_283));
   NAND2_X1 i_1367 (.A1(B[10]), .A2(A[3]), .ZN(n_284));
   AOI22_X1 i_1368 (.A1(B[8]), .A2(A[5]), .B1(B[9]), .B2(A[4]), .ZN(n_285));
   NOR2_X1 i_1369 (.A1(n_176), .A2(n_287), .ZN(n_286));
   NAND2_X1 i_1370 (.A1(B[9]), .A2(A[5]), .ZN(n_287));
   AOI21_X1 i_1371 (.A(n_313), .B1(n_312), .B2(n_305), .ZN(n_304));
   XOR2_X1 i_1372 (.A(n_307), .B(n_306), .Z(n_305));
   NOR2_X1 i_1373 (.A1(n_340), .A2(n_339), .ZN(n_306));
   NOR2_X1 i_1374 (.A1(n_309), .A2(n_308), .ZN(n_307));
   AOI22_X1 i_1375 (.A1(B[3]), .A2(A[10]), .B1(B[2]), .B2(A[11]), .ZN(n_308));
   NOR2_X1 i_1376 (.A1(n_261), .A2(n_311), .ZN(n_309));
   NAND2_X1 i_1377 (.A1(B[3]), .A2(A[11]), .ZN(n_311));
   AOI21_X1 i_1378 (.A(n_313), .B1(n_319), .B2(n_314), .ZN(n_312));
   NOR2_X1 i_1379 (.A1(n_319), .A2(n_314), .ZN(n_313));
   AOI21_X1 i_1380 (.A(n_323), .B1(n_269), .B2(n_321), .ZN(n_314));
   XOR2_X1 i_1381 (.A(n_264), .B(n_320), .Z(n_319));
   NAND2_X1 i_1382 (.A1(n_265), .A2(n_259), .ZN(n_320));
   AOI21_X1 i_1383 (.A(n_323), .B1(n_326), .B2(n_324), .ZN(n_321));
   NOR2_X1 i_1384 (.A1(n_326), .A2(n_324), .ZN(n_323));
   NAND2_X1 i_1385 (.A1(n_330), .A2(n_325), .ZN(n_324));
   NAND2_X1 i_1386 (.A1(n_328), .A2(n_327), .ZN(n_325));
   AOI21_X1 i_1387 (.A(n_335), .B1(n_333), .B2(n_332), .ZN(n_326));
   OR2_X1 i_1388 (.A1(n_272), .A2(n_331), .ZN(n_327));
   NAND2_X1 i_1389 (.A1(B[5]), .A2(A[6]), .ZN(n_328));
   NAND2_X1 i_1390 (.A1(n_272), .A2(n_331), .ZN(n_330));
   NAND2_X1 i_1391 (.A1(B[3]), .A2(A[8]), .ZN(n_331));
   NOR2_X1 i_1392 (.A1(n_339), .A2(n_29), .ZN(n_332));
   NOR2_X1 i_1393 (.A1(n_335), .A2(n_334), .ZN(n_333));
   AOI22_X1 i_1394 (.A1(B[1]), .A2(A[10]), .B1(B[0]), .B2(A[11]), .ZN(n_334));
   NOR2_X1 i_1395 (.A1(n_260), .A2(n_338), .ZN(n_335));
   NAND2_X1 i_1396 (.A1(B[0]), .A2(A[10]), .ZN(n_338));
   INV_X1 i_1397 (.A(A[9]), .ZN(n_339));
   INV_X1 i_1398 (.A(B[4]), .ZN(n_340));
   AOI22_X1 i_1399 (.A1(n_357), .A2(n_356), .B1(n_375), .B2(n_355), .ZN(n_354));
   XOR2_X1 i_1400 (.A(n_357), .B(n_356), .Z(n_355));
   XOR2_X1 i_1401 (.A(n_359), .B(n_358), .Z(n_356));
   XNOR2_X1 i_1402 (.A(n_198), .B(n_371), .ZN(n_357));
   NOR2_X1 i_1403 (.A1(n_425), .A2(n_99), .ZN(n_358));
   NOR2_X1 i_1404 (.A1(n_369), .A2(n_368), .ZN(n_359));
   AOI22_X1 i_1405 (.A1(B[6]), .A2(A[5]), .B1(B[7]), .B2(A[4]), .ZN(n_368));
   NOR2_X1 i_1406 (.A1(n_175), .A2(n_370), .ZN(n_369));
   NAND2_X1 i_1407 (.A1(B[6]), .A2(A[4]), .ZN(n_370));
   NOR2_X1 i_1408 (.A1(n_373), .A2(n_372), .ZN(n_371));
   AOI22_X1 i_1409 (.A1(B[9]), .A2(A[2]), .B1(B[10]), .B2(A[1]), .ZN(n_372));
   NOR2_X1 i_1410 (.A1(n_208), .A2(n_374), .ZN(n_373));
   NAND2_X1 i_1411 (.A1(B[9]), .A2(A[1]), .ZN(n_374));
   OAI22_X1 i_1412 (.A1(n_379), .A2(n_377), .B1(n_390), .B2(n_376), .ZN(n_375));
   XNOR2_X1 i_1413 (.A(n_379), .B(n_377), .ZN(n_376));
   INV_X1 i_1414 (.A(n_378), .ZN(n_377));
   OAI22_X1 i_1415 (.A1(n_396), .A2(n_389), .B1(n_388), .B2(n_387), .ZN(n_378));
   AOI21_X1 i_1416 (.A(n_384), .B1(n_381), .B2(n_380), .ZN(n_379));
   NOR2_X1 i_1417 (.A1(n_426), .A2(n_31), .ZN(n_380));
   NOR2_X1 i_1418 (.A1(n_384), .A2(n_382), .ZN(n_381));
   AOI22_X1 i_1419 (.A1(B[8]), .A2(A[1]), .B1(B[7]), .B2(A[2]), .ZN(n_382));
   NOR2_X1 i_1420 (.A1(n_386), .A2(n_385), .ZN(n_384));
   NAND2_X1 i_1421 (.A1(B[8]), .A2(A[2]), .ZN(n_385));
   NAND2_X1 i_1422 (.A1(B[7]), .A2(A[1]), .ZN(n_386));
   NAND2_X1 i_1423 (.A1(B[6]), .A2(A[3]), .ZN(n_387));
   XNOR2_X1 i_1424 (.A(n_396), .B(n_389), .ZN(n_388));
   NAND2_X1 i_1425 (.A1(B[5]), .A2(A[4]), .ZN(n_389));
   AOI21_X1 i_1426 (.A(n_398), .B1(n_397), .B2(n_391), .ZN(n_390));
   OAI21_X1 i_1427 (.A(n_395), .B1(n_393), .B2(n_392), .ZN(n_391));
   NAND2_X1 i_1428 (.A1(B[5]), .A2(A[3]), .ZN(n_392));
   NAND2_X1 i_1429 (.A1(n_395), .A2(n_394), .ZN(n_393));
   OAI22_X1 i_1430 (.A1(n_424), .A2(n_423), .B1(n_422), .B2(n_340), .ZN(n_394));
   OR3_X1 i_1431 (.A1(n_424), .A2(n_396), .A3(n_422), .ZN(n_395));
   NAND2_X1 i_1432 (.A1(B[4]), .A2(A[5]), .ZN(n_396));
   AOI21_X1 i_1433 (.A(n_398), .B1(n_400), .B2(n_399), .ZN(n_397));
   NOR2_X1 i_1434 (.A1(n_400), .A2(n_399), .ZN(n_398));
   AOI21_X1 i_1435 (.A(n_419), .B1(n_417), .B2(n_416), .ZN(n_399));
   OR2_X1 i_1436 (.A1(n_28), .A2(n_339), .ZN(n_400));
   NOR2_X1 i_1437 (.A1(n_29), .A2(n_170), .ZN(n_416));
   NOR2_X1 i_1438 (.A1(n_419), .A2(n_418), .ZN(n_417));
   AOI22_X1 i_1439 (.A1(B[0]), .A2(A[8]), .B1(B[1]), .B2(A[7]), .ZN(n_418));
   NOR2_X1 i_1440 (.A1(n_421), .A2(n_420), .ZN(n_419));
   NAND2_X1 i_1441 (.A1(B[1]), .A2(A[8]), .ZN(n_420));
   NAND2_X1 i_1442 (.A1(B[0]), .A2(A[7]), .ZN(n_421));
   INV_X1 i_1443 (.A(A[4]), .ZN(n_422));
   INV_X1 i_1444 (.A(A[5]), .ZN(n_423));
   INV_X1 i_1445 (.A(B[3]), .ZN(n_424));
   INV_X1 i_1446 (.A(B[8]), .ZN(n_425));
   INV_X1 i_1447 (.A(B[9]), .ZN(n_426));
   AOI21_X1 i_1448 (.A(n_441), .B1(n_439), .B2(n_437), .ZN(n_427));
   XOR2_X1 i_1449 (.A(n_328), .B(n_438), .Z(n_437));
   NAND2_X1 i_1450 (.A1(n_327), .A2(n_330), .ZN(n_438));
   AOI21_X1 i_1451 (.A(n_441), .B1(n_444), .B2(n_442), .ZN(n_439));
   NOR2_X1 i_1452 (.A1(n_444), .A2(n_442), .ZN(n_441));
   XNOR2_X1 i_1453 (.A(n_333), .B(n_332), .ZN(n_442));
   AOI22_X1 i_1454 (.A1(n_457), .A2(n_453), .B1(n_446), .B2(n_445), .ZN(n_444));
   NOR2_X1 i_1455 (.A1(n_257), .A2(n_339), .ZN(n_445));
   XOR2_X1 i_1456 (.A(n_457), .B(n_453), .Z(n_446));
   OAI33_X1 i_1457 (.A1(n_424), .A2(n_170), .A3(n_454), .B1(n_458), .B2(n_257), 
      .B3(n_455), .ZN(n_453));
   XNOR2_X1 i_1458 (.A(n_420), .B(n_455), .ZN(n_454));
   NAND2_X1 i_1459 (.A1(B[2]), .A2(A[7]), .ZN(n_455));
   INV_X1 i_1460 (.A(n_338), .ZN(n_457));
   INV_X1 i_1461 (.A(A[8]), .ZN(n_458));
   INV_X1 i_1462 (.A(n_460), .ZN(n_459));
   OAI21_X1 i_1463 (.A(n_496), .B1(n_495), .B2(n_461), .ZN(n_460));
   AOI22_X1 i_1464 (.A1(n_488), .A2(n_487), .B1(n_470), .B2(n_462), .ZN(n_461));
   OAI21_X1 i_1465 (.A(n_468), .B1(n_466), .B2(n_465), .ZN(n_462));
   NAND2_X1 i_1466 (.A1(B[2]), .A2(A[12]), .ZN(n_465));
   NAND2_X1 i_1467 (.A1(n_468), .A2(n_467), .ZN(n_466));
   OAI22_X1 i_1468 (.A1(n_557), .A2(n_28), .B1(n_256), .B2(n_257), .ZN(n_467));
   OR3_X1 i_1469 (.A1(n_28), .A2(n_469), .A3(n_256), .ZN(n_468));
   NAND2_X1 i_1470 (.A1(B[1]), .A2(A[14]), .ZN(n_469));
   XOR2_X1 i_1471 (.A(n_488), .B(n_487), .Z(n_470));
   OAI22_X1 i_1472 (.A1(n_311), .A2(n_494), .B1(n_492), .B2(n_489), .ZN(n_487));
   NOR2_X1 i_1473 (.A1(n_558), .A2(n_28), .ZN(n_488));
   NAND2_X1 i_1474 (.A1(B[5]), .A2(A[9]), .ZN(n_489));
   XNOR2_X1 i_1475 (.A(n_311), .B(n_494), .ZN(n_492));
   NAND2_X1 i_1476 (.A1(B[4]), .A2(A[10]), .ZN(n_494));
   OAI21_X1 i_1477 (.A(n_496), .B1(n_501), .B2(n_498), .ZN(n_495));
   NAND2_X1 i_1478 (.A1(n_501), .A2(n_498), .ZN(n_496));
   OAI22_X1 i_1479 (.A1(n_533), .A2(n_532), .B1(n_530), .B2(n_516), .ZN(n_498));
   OAI33_X1 i_1480 (.A1(n_560), .A2(n_31), .A3(n_502), .B1(n_33), .B2(n_229), 
      .B3(n_515), .ZN(n_501));
   XNOR2_X1 i_1481 (.A(n_521), .B(n_515), .ZN(n_502));
   NAND2_X1 i_1482 (.A1(B[14]), .A2(A[1]), .ZN(n_515));
   OAI21_X1 i_1483 (.A(n_522), .B1(n_520), .B2(n_517), .ZN(n_516));
   NOR2_X1 i_1484 (.A1(n_559), .A2(n_31), .ZN(n_517));
   NOR2_X1 i_1485 (.A1(n_204), .A2(n_521), .ZN(n_520));
   NAND2_X1 i_1486 (.A1(B[13]), .A2(A[2]), .ZN(n_521));
   INV_X1 i_1487 (.A(n_523), .ZN(n_522));
   AOI22_X1 i_1488 (.A1(B[12]), .A2(A[2]), .B1(B[13]), .B2(A[1]), .ZN(n_523));
   OAI21_X1 i_1489 (.A(n_531), .B1(n_533), .B2(n_532), .ZN(n_524));
   INV_X1 i_1490 (.A(n_531), .ZN(n_530));
   NAND2_X1 i_1491 (.A1(n_533), .A2(n_532), .ZN(n_531));
   OAI21_X1 i_1492 (.A(n_536), .B1(n_555), .B2(n_534), .ZN(n_532));
   AOI21_X1 i_1493 (.A(n_543), .B1(n_541), .B2(n_540), .ZN(n_533));
   NOR2_X1 i_1494 (.A1(n_284), .A2(n_535), .ZN(n_534));
   NAND2_X1 i_1495 (.A1(B[11]), .A2(A[4]), .ZN(n_535));
   INV_X1 i_1496 (.A(n_537), .ZN(n_536));
   AOI22_X1 i_1497 (.A1(B[11]), .A2(A[3]), .B1(B[10]), .B2(A[4]), .ZN(n_537));
   NOR2_X1 i_1498 (.A1(n_170), .A2(n_425), .ZN(n_540));
   NOR2_X1 i_1499 (.A1(n_543), .A2(n_542), .ZN(n_541));
   AOI22_X1 i_1500 (.A1(B[7]), .A2(A[7]), .B1(B[6]), .B2(A[8]), .ZN(n_542));
   NOR3_X1 i_1501 (.A1(n_169), .A2(n_544), .A3(n_556), .ZN(n_543));
   NAND2_X1 i_1502 (.A1(B[7]), .A2(A[8]), .ZN(n_544));
   INV_X1 i_1503 (.A(n_287), .ZN(n_555));
   INV_X1 i_1504 (.A(A[7]), .ZN(n_556));
   INV_X1 i_1505 (.A(A[14]), .ZN(n_557));
   INV_X1 i_1506 (.A(A[15]), .ZN(n_558));
   INV_X1 i_1507 (.A(B[14]), .ZN(n_559));
   INV_X1 i_1508 (.A(B[15]), .ZN(n_560));
   NAND2_X1 i_1509 (.A1(B[5]), .A2(A[11]), .ZN(n_561));
   NOR2_X1 i_1510 (.A1(n_561), .A2(n_494), .ZN(n_562));
   AOI22_X1 i_1511 (.A1(B[5]), .A2(A[10]), .B1(B[4]), .B2(A[11]), .ZN(n_564));
   NOR2_X1 i_1512 (.A1(n_562), .A2(n_564), .ZN(n_565));
   NOR2_X1 i_1513 (.A1(n_169), .A2(n_339), .ZN(n_566));
   NAND2_X1 i_1514 (.A1(B[8]), .A2(A[7]), .ZN(n_567));
   NAND2_X1 i_1515 (.A1(n_567), .A2(n_544), .ZN(n_568));
   NAND2_X1 i_1516 (.A1(B[9]), .A2(A[6]), .ZN(n_569));
   NOR2_X1 i_1517 (.A1(n_567), .A2(n_544), .ZN(n_570));
   INV_X1 i_1518 (.A(n_570), .ZN(n_571));
   AOI21_X1 i_1519 (.A(n_562), .B1(n_565), .B2(n_566), .ZN(n_572));
   INV_X1 i_1520 (.A(n_569), .ZN(n_573));
   OAI21_X1 i_1521 (.A(n_568), .B1(n_570), .B2(n_573), .ZN(n_574));
   NOR2_X1 i_1522 (.A1(n_572), .A2(n_574), .ZN(n_575));
   AOI21_X1 i_1523 (.A(n_575), .B1(n_572), .B2(n_574), .ZN(n_576));
   INV_X1 i_1524 (.A(n_535), .ZN(n_577));
   AOI21_X1 i_1525 (.A(n_577), .B1(B[12]), .B2(A[3]), .ZN(n_578));
   NAND2_X1 i_1526 (.A1(B[10]), .A2(A[5]), .ZN(n_579));
   NAND3_X1 i_1527 (.A1(n_577), .A2(B[12]), .A3(A[3]), .ZN(n_580));
   AOI21_X1 i_1528 (.A(n_578), .B1(n_579), .B2(n_580), .ZN(n_581));
   AOI21_X1 i_1529 (.A(n_575), .B1(n_576), .B2(n_581), .ZN(n_582));
   NAND2_X1 i_1530 (.A1(B[15]), .A2(A[2]), .ZN(n_583));
   NOR2_X1 i_1531 (.A1(n_583), .A2(n_515), .ZN(n_589));
   AOI22_X1 i_1532 (.A1(B[15]), .A2(A[1]), .B1(B[14]), .B2(A[2]), .ZN(n_590));
   NOR2_X1 i_1533 (.A1(n_589), .A2(n_590), .ZN(n_591));
   INV_X1 i_1534 (.A(B[16]), .ZN(n_592));
   NOR2_X1 i_1535 (.A1(n_592), .A2(n_31), .ZN(n_593));
   AOI21_X1 i_1536 (.A(n_589), .B1(n_591), .B2(n_593), .ZN(n_598));
   NAND2_X1 i_1537 (.A1(B[12]), .A2(A[5]), .ZN(n_599));
   AOI22_X1 i_1538 (.A1(B[12]), .A2(A[4]), .B1(B[11]), .B2(A[5]), .ZN(n_600));
   NAND2_X1 i_1539 (.A1(B[13]), .A2(A[3]), .ZN(n_601));
   NOR2_X1 i_1540 (.A1(n_599), .A2(n_535), .ZN(n_602));
   INV_X1 i_1541 (.A(n_602), .ZN(n_603));
   OAI21_X1 i_1542 (.A(n_603), .B1(n_600), .B2(n_601), .ZN(n_604));
   XNOR2_X1 i_1543 (.A(n_598), .B(n_604), .ZN(n_605));
   XOR2_X1 i_1544 (.A(n_582), .B(n_605), .Z(n_606));
   NAND2_X1 i_1545 (.A1(B[16]), .A2(A[1]), .ZN(n_607));
   XNOR2_X1 i_1546 (.A(n_583), .B(n_607), .ZN(n_608));
   NAND2_X1 i_1547 (.A1(B[17]), .A2(A[0]), .ZN(n_609));
   XNOR2_X1 i_1548 (.A(n_608), .B(n_609), .ZN(n_610));
   XOR2_X1 i_1549 (.A(n_606), .B(n_610), .Z(n_611));
   NAND2_X1 i_1550 (.A1(A[16]), .A2(B[1]), .ZN(n_612));
   NAND2_X1 i_1551 (.A1(A[13]), .A2(B[2]), .ZN(n_613));
   XNOR2_X1 i_1552 (.A(n_613), .B(n_469), .ZN(n_614));
   NAND2_X1 i_1553 (.A1(A[12]), .A2(B[3]), .ZN(n_615));
   NAND2_X1 i_1554 (.A1(B[0]), .A2(A[17]), .ZN(n_616));
   XNOR2_X1 i_1555 (.A(n_612), .B(n_616), .ZN(n_640));
   NAND2_X1 i_1556 (.A1(A[15]), .A2(B[2]), .ZN(n_645));
   AOI22_X1 i_1557 (.A1(B[0]), .A2(A[16]), .B1(A[15]), .B2(B[1]), .ZN(n_647));
   INV_X1 i_1558 (.A(n_647), .ZN(n_660));
   OAI22_X1 i_1559 (.A1(n_614), .A2(n_615), .B1(n_613), .B2(n_469), .ZN(n_661));
   INV_X1 i_1560 (.A(n_488), .ZN(n_662));
   NOR2_X1 i_1561 (.A1(n_612), .A2(n_662), .ZN(n_663));
   OAI21_X1 i_1562 (.A(n_660), .B1(n_661), .B2(n_663), .ZN(n_664));
   XNOR2_X1 i_1563 (.A(n_640), .B(n_645), .ZN(n_665));
   XNOR2_X1 i_1564 (.A(n_664), .B(n_665), .ZN(n_666));
   NAND2_X1 i_1565 (.A1(B[3]), .A2(A[14]), .ZN(n_667));
   NAND2_X1 i_1566 (.A1(B[4]), .A2(A[13]), .ZN(n_668));
   XNOR2_X1 i_1567 (.A(n_667), .B(n_668), .ZN(n_669));
   NAND2_X1 i_1568 (.A1(A[12]), .A2(B[5]), .ZN(n_670));
   XNOR2_X1 i_1569 (.A(n_669), .B(n_670), .ZN(n_671));
   NAND2_X1 i_1570 (.A1(A[10]), .A2(B[6]), .ZN(n_675));
   XNOR2_X1 i_1571 (.A(n_675), .B(n_561), .ZN(n_676));
   NAND2_X1 i_1572 (.A1(A[9]), .A2(B[7]), .ZN(n_677));
   OAI22_X1 i_1573 (.A1(n_676), .A2(n_677), .B1(n_675), .B2(n_561), .ZN(n_678));
   NOR2_X1 i_1574 (.A1(n_613), .A2(n_667), .ZN(n_679));
   INV_X1 i_1575 (.A(n_679), .ZN(n_680));
   AOI22_X1 i_1576 (.A1(A[13]), .A2(B[3]), .B1(A[14]), .B2(B[2]), .ZN(n_681));
   OR2_X1 i_1577 (.A1(n_679), .A2(n_681), .ZN(n_682));
   OR2_X1 i_1578 (.A1(n_340), .A2(n_258), .ZN(n_683));
   OAI21_X1 i_1579 (.A(n_680), .B1(n_682), .B2(n_683), .ZN(n_684));
   NAND2_X1 i_1580 (.A1(n_678), .A2(n_684), .ZN(n_685));
   OAI21_X1 i_1581 (.A(n_685), .B1(n_678), .B2(n_684), .ZN(n_686));
   AOI22_X1 i_1582 (.A1(A[7]), .A2(B[9]), .B1(A[8]), .B2(B[8]), .ZN(n_687));
   INV_X1 i_1583 (.A(n_687), .ZN(n_689));
   NOR3_X1 i_1584 (.A1(n_567), .A2(n_426), .A3(n_458), .ZN(n_690));
   AND2_X1 i_1585 (.A1(A[6]), .A2(B[10]), .ZN(n_691));
   OAI21_X1 i_1586 (.A(n_689), .B1(n_690), .B2(n_691), .ZN(n_692));
   OAI21_X1 i_1587 (.A(n_685), .B1(n_686), .B2(n_692), .ZN(n_693));
   INV_X1 i_1588 (.A(n_693), .ZN(n_694));
   NAND2_X1 i_1589 (.A1(B[2]), .A2(A[17]), .ZN(n_695));
   NOR2_X1 i_1590 (.A1(n_612), .A2(n_695), .ZN(n_696));
   AOI22_X1 i_1591 (.A1(A[16]), .A2(B[2]), .B1(A[17]), .B2(B[1]), .ZN(n_726));
   NOR2_X1 i_1592 (.A1(n_696), .A2(n_726), .ZN(n_731));
   NOR2_X1 i_1593 (.A1(n_424), .A2(n_558), .ZN(n_737));
   OAI22_X1 i_1594 (.A1(n_608), .A2(n_609), .B1(n_583), .B2(n_607), .ZN(n_750));
   XNOR2_X1 i_1595 (.A(n_731), .B(n_737), .ZN(n_760));
   XOR2_X1 i_1596 (.A(n_760), .B(n_750), .Z(n_761));
   NOR2_X1 i_1597 (.A1(n_687), .A2(n_690), .ZN(n_762));
   XNOR2_X1 i_1598 (.A(n_762), .B(n_691), .ZN(n_763));
   NOR2_X1 i_1599 (.A1(n_602), .A2(n_600), .ZN(n_769));
   XOR2_X1 i_1600 (.A(n_769), .B(n_601), .Z(n_770));
   NOR2_X1 i_1601 (.A1(n_763), .A2(n_770), .ZN(n_771));
   AOI21_X1 i_1602 (.A(n_771), .B1(n_770), .B2(n_763), .ZN(n_772));
   XOR2_X1 i_1603 (.A(n_591), .B(n_593), .Z(n_773));
   AOI21_X1 i_1604 (.A(n_771), .B1(n_772), .B2(n_773), .ZN(n_774));
   XNOR2_X1 i_1605 (.A(n_686), .B(n_692), .ZN(n_775));
   NOR2_X1 i_1606 (.A1(n_774), .A2(n_775), .ZN(n_776));
   AOI21_X1 i_1607 (.A(n_776), .B1(n_774), .B2(n_775), .ZN(n_777));
   NOR2_X1 i_1608 (.A1(n_663), .A2(n_647), .ZN(n_778));
   XOR2_X1 i_1609 (.A(n_661), .B(n_778), .Z(n_779));
   XOR2_X1 i_1610 (.A(n_682), .B(n_683), .Z(n_780));
   XOR2_X1 i_1611 (.A(n_779), .B(n_780), .Z(n_781));
   XOR2_X1 i_1612 (.A(n_676), .B(n_677), .Z(n_782));
   AOI22_X1 i_1613 (.A1(n_781), .A2(n_782), .B1(n_779), .B2(n_780), .ZN(n_783));
   INV_X1 i_1614 (.A(n_783), .ZN(n_784));
   AOI21_X1 i_1615 (.A(n_776), .B1(n_777), .B2(n_784), .ZN(n_802));
   XNOR2_X1 i_1616 (.A(n_693), .B(n_761), .ZN(n_817));
   OAI22_X1 i_1617 (.A1(n_666), .A2(n_671), .B1(n_664), .B2(n_665), .ZN(n_829));
   NAND2_X1 i_1618 (.A1(n_817), .A2(n_829), .ZN(n_830));
   OAI21_X1 i_1619 (.A(n_830), .B1(n_829), .B2(n_817), .ZN(n_831));
   OAI21_X1 i_1620 (.A(n_830), .B1(n_802), .B2(n_831), .ZN(n_832));
   XNOR2_X1 i_1621 (.A(n_840), .B(n_834), .ZN(n_833));
   XOR2_X1 i_1622 (.A(n_836), .B(n_835), .Z(n_834));
   NAND2_X1 i_1623 (.A1(n_838), .A2(n_837), .ZN(n_835));
   NAND2_X1 i_1624 (.A1(B[4]), .A2(A[15]), .ZN(n_836));
   NAND2_X1 i_1625 (.A1(n_695), .A2(n_839), .ZN(n_837));
   OR2_X1 i_1626 (.A1(n_695), .A2(n_839), .ZN(n_838));
   NAND2_X1 i_1627 (.A1(B[3]), .A2(A[16]), .ZN(n_839));
   XOR2_X1 i_1628 (.A(n_847), .B(n_841), .Z(n_840));
   XNOR2_X1 i_1629 (.A(n_846), .B(n_842), .ZN(n_841));
   NOR2_X1 i_1630 (.A1(n_845), .A2(n_843), .ZN(n_842));
   AOI22_X1 i_1631 (.A1(B[0]), .A2(A[19]), .B1(B[1]), .B2(A[18]), .ZN(n_843));
   INV_X1 i_1632 (.A(n_845), .ZN(n_844));
   NOR3_X1 i_1633 (.A1(n_257), .A2(n_848), .A3(n_853), .ZN(n_845));
   AOI21_X1 i_1634 (.A(n_696), .B1(n_731), .B2(n_737), .ZN(n_846));
   OAI21_X1 i_1635 (.A(n_850), .B1(n_849), .B2(n_848), .ZN(n_847));
   NAND2_X1 i_1636 (.A1(B[0]), .A2(A[18]), .ZN(n_848));
   OAI21_X1 i_1637 (.A(n_850), .B1(n_852), .B2(n_851), .ZN(n_849));
   NAND2_X1 i_1638 (.A1(n_852), .A2(n_851), .ZN(n_850));
   OAI22_X1 i_1639 (.A1(n_667), .A2(n_668), .B1(n_669), .B2(n_670), .ZN(n_851));
   OAI22_X1 i_1640 (.A1(n_612), .A2(n_616), .B1(n_640), .B2(n_645), .ZN(n_852));
   INV_X1 i_1641 (.A(A[19]), .ZN(n_853));
   NAND2_X1 i_1642 (.A1(B[19]), .A2(A[2]), .ZN(n_855));
   INV_X1 i_1643 (.A(B[20]), .ZN(n_856));
   NOR2_X1 i_1644 (.A1(n_856), .A2(n_31), .ZN(n_857));
   NAND3_X1 i_1645 (.A1(n_857), .A2(A[1]), .A3(B[21]), .ZN(n_860));
   AOI22_X1 i_1646 (.A1(B[20]), .A2(A[1]), .B1(B[21]), .B2(A[0]), .ZN(n_884));
   INV_X1 i_1647 (.A(n_860), .ZN(n_885));
   NOR2_X1 i_1648 (.A1(n_885), .A2(n_884), .ZN(n_886));
   XNOR2_X1 i_1649 (.A(n_886), .B(n_855), .ZN(n_887));
   NAND2_X1 i_1650 (.A1(B[18]), .A2(A[3]), .ZN(n_888));
   NAND2_X1 i_1651 (.A1(A[5]), .A2(B[17]), .ZN(n_889));
   AOI22_X1 i_1652 (.A1(B[16]), .A2(A[5]), .B1(B[17]), .B2(A[4]), .ZN(n_896));
   NOR3_X1 i_1653 (.A1(n_889), .A2(n_422), .A3(n_592), .ZN(n_897));
   NOR2_X1 i_1654 (.A1(n_897), .A2(n_896), .ZN(n_898));
   XNOR2_X1 i_1655 (.A(n_898), .B(n_888), .ZN(n_899));
   XOR2_X1 i_1656 (.A(n_899), .B(n_887), .Z(n_901));
   INV_X1 i_1657 (.A(n_897), .ZN(n_902));
   XOR2_X1 i_1658 (.A(n_944), .B(n_904), .Z(n_903));
   AOI22_X1 i_1659 (.A1(n_943), .A2(n_941), .B1(n_940), .B2(n_905), .ZN(n_904));
   AOI22_X1 i_1660 (.A1(n_927), .A2(n_925), .B1(n_924), .B2(n_906), .ZN(n_905));
   OAI21_X1 i_1661 (.A(n_909), .B1(n_857), .B2(n_910), .ZN(n_906));
   NAND2_X1 i_1662 (.A1(n_857), .A2(n_910), .ZN(n_909));
   NOR2_X1 i_1663 (.A1(n_912), .A2(n_911), .ZN(n_910));
   AOI22_X1 i_1664 (.A1(B[18]), .A2(A[2]), .B1(B[19]), .B2(A[1]), .ZN(n_911));
   NOR2_X1 i_1665 (.A1(n_855), .A2(n_913), .ZN(n_912));
   NAND2_X1 i_1666 (.A1(B[18]), .A2(A[1]), .ZN(n_913));
   XOR2_X1 i_1667 (.A(n_927), .B(n_925), .Z(n_924));
   XOR2_X1 i_1668 (.A(n_929), .B(n_926), .Z(n_925));
   NAND2_X1 i_1669 (.A1(B[17]), .A2(A[3]), .ZN(n_926));
   XNOR2_X1 i_1670 (.A(n_1003), .B(n_1002), .ZN(n_927));
   INV_X1 i_1671 (.A(n_929), .ZN(n_928));
   XOR2_X1 i_1672 (.A(n_939), .B(n_938), .Z(n_929));
   NAND2_X1 i_1673 (.A1(B[15]), .A2(A[5]), .ZN(n_938));
   NAND2_X1 i_1674 (.A1(B[16]), .A2(A[4]), .ZN(n_939));
   XOR2_X1 i_1675 (.A(n_943), .B(n_941), .Z(n_940));
   XOR2_X1 i_1676 (.A(n_988), .B(n_942), .Z(n_941));
   OAI21_X1 i_1677 (.A(n_985), .B1(n_987), .B2(n_986), .ZN(n_942));
   XOR2_X1 i_1678 (.A(n_1001), .B(n_1000), .Z(n_943));
   XNOR2_X1 i_1679 (.A(n_955), .B(n_945), .ZN(n_944));
   XOR2_X1 i_1680 (.A(n_950), .B(n_946), .Z(n_945));
   OR2_X1 i_1681 (.A1(n_948), .A2(n_947), .ZN(n_946));
   AOI22_X1 i_1682 (.A1(B[0]), .A2(A[22]), .B1(B[1]), .B2(A[21]), .ZN(n_947));
   NOR2_X1 i_1683 (.A1(n_988), .A2(n_949), .ZN(n_948));
   NAND2_X1 i_1684 (.A1(B[1]), .A2(A[22]), .ZN(n_949));
   OAI21_X1 i_1685 (.A(n_953), .B1(n_952), .B2(n_951), .ZN(n_950));
   NOR2_X1 i_1686 (.A1(n_1028), .A2(n_424), .ZN(n_951));
   NOR2_X1 i_1687 (.A1(n_993), .A2(n_954), .ZN(n_952));
   NAND2_X1 i_1688 (.A1(n_993), .A2(n_954), .ZN(n_953));
   NAND2_X1 i_1689 (.A1(B[2]), .A2(A[19]), .ZN(n_954));
   XNOR2_X1 i_1690 (.A(n_999), .B(n_978), .ZN(n_955));
   OAI22_X1 i_1691 (.A1(n_987), .A2(n_986), .B1(n_988), .B2(n_984), .ZN(n_978));
   INV_X1 i_1692 (.A(n_985), .ZN(n_984));
   NAND2_X1 i_1693 (.A1(n_987), .A2(n_986), .ZN(n_985));
   AOI21_X1 i_1694 (.A(n_992), .B1(n_990), .B2(n_989), .ZN(n_986));
   AOI21_X1 i_1695 (.A(n_998), .B1(n_995), .B2(n_994), .ZN(n_987));
   NAND2_X1 i_1696 (.A1(B[0]), .A2(A[21]), .ZN(n_988));
   NOR2_X1 i_1697 (.A1(n_1028), .A2(n_29), .ZN(n_989));
   NOR2_X1 i_1698 (.A1(n_992), .A2(n_991), .ZN(n_990));
   AOI22_X1 i_1699 (.A1(B[0]), .A2(A[20]), .B1(B[1]), .B2(A[19]), .ZN(n_991));
   NOR3_X1 i_1700 (.A1(n_28), .A2(n_993), .A3(n_853), .ZN(n_992));
   NAND2_X1 i_1701 (.A1(B[1]), .A2(A[20]), .ZN(n_993));
   NOR2_X1 i_1702 (.A1(n_1029), .A2(n_558), .ZN(n_994));
   NOR2_X1 i_1703 (.A1(n_998), .A2(n_996), .ZN(n_995));
   AOI22_X1 i_1704 (.A1(B[3]), .A2(A[17]), .B1(B[4]), .B2(A[16]), .ZN(n_996));
   NOR3_X1 i_1705 (.A1(n_839), .A2(n_340), .A3(n_1027), .ZN(n_998));
   AOI21_X1 i_1706 (.A(n_1004), .B1(n_1001), .B2(n_1000), .ZN(n_999));
   AOI21_X1 i_1707 (.A(n_1004), .B1(n_1006), .B2(n_1005), .ZN(n_1000));
   OAI22_X1 i_1708 (.A1(n_1008), .A2(n_1007), .B1(n_1003), .B2(n_1002), .ZN(
      n_1001));
   NAND2_X1 i_1709 (.A1(B[14]), .A2(A[6]), .ZN(n_1002));
   XNOR2_X1 i_1710 (.A(n_1008), .B(n_1007), .ZN(n_1003));
   NOR2_X1 i_1711 (.A1(n_1006), .A2(n_1005), .ZN(n_1004));
   AOI21_X1 i_1712 (.A(n_1015), .B1(n_1013), .B2(n_1009), .ZN(n_1005));
   AOI21_X1 i_1713 (.A(n_1024), .B1(n_1022), .B2(n_1018), .ZN(n_1006));
   NAND2_X1 i_1714 (.A1(B[13]), .A2(A[7]), .ZN(n_1007));
   NAND2_X1 i_1715 (.A1(B[12]), .A2(A[8]), .ZN(n_1008));
   INV_X1 i_1716 (.A(n_1011), .ZN(n_1009));
   NAND2_X1 i_1717 (.A1(B[6]), .A2(A[14]), .ZN(n_1011));
   NOR2_X1 i_1718 (.A1(n_1015), .A2(n_1014), .ZN(n_1013));
   AOI22_X1 i_1719 (.A1(B[8]), .A2(A[12]), .B1(B[7]), .B2(A[13]), .ZN(n_1014));
   NOR2_X1 i_1720 (.A1(n_1017), .A2(n_1016), .ZN(n_1015));
   NAND2_X1 i_1721 (.A1(B[8]), .A2(A[13]), .ZN(n_1016));
   NAND2_X1 i_1722 (.A1(B[7]), .A2(A[12]), .ZN(n_1017));
   INV_X1 i_1723 (.A(n_1021), .ZN(n_1018));
   NAND2_X1 i_1724 (.A1(B[11]), .A2(A[9]), .ZN(n_1021));
   NOR2_X1 i_1725 (.A1(n_1024), .A2(n_1023), .ZN(n_1022));
   AOI22_X1 i_1726 (.A1(B[9]), .A2(A[11]), .B1(B[10]), .B2(A[10]), .ZN(n_1023));
   NOR2_X1 i_1727 (.A1(n_1026), .A2(n_1025), .ZN(n_1024));
   NAND2_X1 i_1728 (.A1(B[10]), .A2(A[11]), .ZN(n_1025));
   NAND2_X1 i_1729 (.A1(B[9]), .A2(A[10]), .ZN(n_1026));
   INV_X1 i_1730 (.A(A[17]), .ZN(n_1027));
   INV_X1 i_1731 (.A(A[18]), .ZN(n_1028));
   INV_X1 i_1732 (.A(B[5]), .ZN(n_1029));
   INV_X1 i_1733 (.A(n_1031), .ZN(n_1030));
   AOI22_X1 i_1734 (.A1(n_1034), .A2(n_1033), .B1(n_1096), .B2(n_1032), .ZN(
      n_1031));
   XOR2_X1 i_1735 (.A(n_1034), .B(n_1033), .Z(n_1032));
   XNOR2_X1 i_1736 (.A(n_1061), .B(n_1056), .ZN(n_1033));
   OAI21_X1 i_1737 (.A(n_1053), .B1(n_1052), .B2(n_1035), .ZN(n_1034));
   XOR2_X1 i_1738 (.A(n_1048), .B(n_1036), .Z(n_1035));
   NOR2_X1 i_1739 (.A1(n_170), .A2(n_560), .ZN(n_1036));
   NOR2_X1 i_1740 (.A1(n_1050), .A2(n_1049), .ZN(n_1048));
   AOI22_X1 i_1741 (.A1(B[13]), .A2(A[8]), .B1(B[14]), .B2(A[7]), .ZN(n_1049));
   NOR2_X1 i_1742 (.A1(n_1007), .A2(n_1051), .ZN(n_1050));
   NAND2_X1 i_1743 (.A1(B[14]), .A2(A[8]), .ZN(n_1051));
   NOR2_X1 i_1744 (.A1(n_1055), .A2(n_1054), .ZN(n_1052));
   NAND2_X1 i_1745 (.A1(n_1055), .A2(n_1054), .ZN(n_1053));
   XNOR2_X1 i_1746 (.A(n_1025), .B(n_1057), .ZN(n_1054));
   XNOR2_X1 i_1747 (.A(n_1065), .B(n_1064), .ZN(n_1055));
   OAI22_X1 i_1748 (.A1(n_1021), .A2(n_1060), .B1(n_1025), .B2(n_1057), .ZN(
      n_1056));
   OAI21_X1 i_1749 (.A(n_1058), .B1(n_1021), .B2(n_1060), .ZN(n_1057));
   INV_X1 i_1750 (.A(n_1059), .ZN(n_1058));
   AOI22_X1 i_1751 (.A1(B[12]), .A2(A[9]), .B1(B[11]), .B2(A[10]), .ZN(n_1059));
   NAND2_X1 i_1752 (.A1(B[12]), .A2(A[10]), .ZN(n_1060));
   XOR2_X1 i_1753 (.A(n_1063), .B(n_1062), .Z(n_1061));
   OAI22_X1 i_1754 (.A1(n_1102), .A2(n_1101), .B1(n_1100), .B2(n_1098), .ZN(
      n_1062));
   OAI22_X1 i_1755 (.A1(n_1016), .A2(n_1095), .B1(n_1065), .B2(n_1064), .ZN(
      n_1063));
   NAND2_X1 i_1756 (.A1(B[9]), .A2(A[12]), .ZN(n_1064));
   XNOR2_X1 i_1757 (.A(n_1016), .B(n_1095), .ZN(n_1065));
   NAND2_X1 i_1758 (.A1(B[7]), .A2(A[14]), .ZN(n_1095));
   AOI22_X1 i_1759 (.A1(n_1111), .A2(n_1104), .B1(n_1103), .B2(n_1097), .ZN(
      n_1096));
   XNOR2_X1 i_1760 (.A(n_1099), .B(n_1098), .ZN(n_1097));
   NAND2_X1 i_1761 (.A1(B[6]), .A2(A[15]), .ZN(n_1098));
   XOR2_X1 i_1762 (.A(n_1102), .B(n_1101), .Z(n_1099));
   AND2_X1 i_1763 (.A1(n_1102), .A2(n_1101), .ZN(n_1100));
   NAND2_X1 i_1764 (.A1(B[5]), .A2(A[16]), .ZN(n_1101));
   NAND2_X1 i_1765 (.A1(B[4]), .A2(A[17]), .ZN(n_1102));
   XOR2_X1 i_1766 (.A(n_1111), .B(n_1104), .Z(n_1103));
   INV_X1 i_1767 (.A(n_1110), .ZN(n_1104));
   AOI22_X1 i_1768 (.A1(n_1119), .A2(n_1118), .B1(n_1117), .B2(n_1113), .ZN(
      n_1110));
   XOR2_X1 i_1769 (.A(n_951), .B(n_1112), .Z(n_1111));
   NOR2_X1 i_1770 (.A1(n_952), .A2(n_1129), .ZN(n_1112));
   OAI22_X1 i_1771 (.A1(n_1026), .A2(n_1116), .B1(n_1115), .B2(n_1114), .ZN(
      n_1113));
   NAND2_X1 i_1772 (.A1(B[10]), .A2(A[9]), .ZN(n_1114));
   XNOR2_X1 i_1773 (.A(n_1026), .B(n_1116), .ZN(n_1115));
   NAND2_X1 i_1774 (.A1(B[8]), .A2(A[11]), .ZN(n_1116));
   XOR2_X1 i_1775 (.A(n_1119), .B(n_1118), .Z(n_1117));
   AOI21_X1 i_1776 (.A(n_1143), .B1(n_836), .B2(n_838), .ZN(n_1118));
   OAI22_X1 i_1777 (.A1(n_1011), .A2(n_1128), .B1(n_1017), .B2(n_1121), .ZN(
      n_1119));
   NOR2_X1 i_1778 (.A1(n_1122), .A2(n_1121), .ZN(n_1120));
   AOI22_X1 i_1779 (.A1(B[5]), .A2(A[14]), .B1(B[6]), .B2(A[13]), .ZN(n_1121));
   NOR2_X1 i_1780 (.A1(n_1011), .A2(n_1128), .ZN(n_1122));
   NAND2_X1 i_1781 (.A1(B[5]), .A2(A[13]), .ZN(n_1128));
   INV_X1 i_1782 (.A(n_953), .ZN(n_1129));
   INV_X1 i_1783 (.A(n_837), .ZN(n_1143));
   AOI22_X1 i_1784 (.A1(n_1197), .A2(n_1146), .B1(n_1196), .B2(n_1145), .ZN(
      n_1144));
   INV_X1 i_1785 (.A(n_1146), .ZN(n_1145));
   XOR2_X1 i_1786 (.A(n_1153), .B(n_1147), .Z(n_1146));
   OAI22_X1 i_1787 (.A1(n_1152), .A2(n_1151), .B1(n_1150), .B2(n_1148), .ZN(
      n_1147));
   NAND2_X1 i_1788 (.A1(A[15]), .A2(B[8]), .ZN(n_1148));
   XNOR2_X1 i_1789 (.A(n_1152), .B(n_1151), .ZN(n_1150));
   NAND2_X1 i_1790 (.A1(A[16]), .A2(B[7]), .ZN(n_1151));
   NAND2_X1 i_1791 (.A1(A[17]), .A2(B[6]), .ZN(n_1152));
   XOR2_X1 i_1792 (.A(n_1190), .B(n_1154), .Z(n_1153));
   AOI21_X1 i_1793 (.A(n_1159), .B1(n_1160), .B2(n_1157), .ZN(n_1154));
   NAND2_X1 i_1794 (.A1(A[14]), .A2(B[9]), .ZN(n_1157));
   NOR2_X1 i_1795 (.A1(n_1161), .A2(n_1159), .ZN(n_1158));
   AOI22_X1 i_1796 (.A1(A[12]), .A2(B[11]), .B1(A[13]), .B2(B[10]), .ZN(n_1159));
   INV_X1 i_1797 (.A(n_1161), .ZN(n_1160));
   NOR2_X1 i_1798 (.A1(n_1173), .A2(n_1164), .ZN(n_1161));
   NAND2_X1 i_1799 (.A1(A[13]), .A2(B[11]), .ZN(n_1164));
   NAND2_X1 i_1800 (.A1(A[12]), .A2(B[10]), .ZN(n_1173));
   OAI22_X1 i_1801 (.A1(n_1194), .A2(n_1193), .B1(n_1192), .B2(n_1191), .ZN(
      n_1190));
   NAND2_X1 i_1802 (.A1(A[18]), .A2(B[5]), .ZN(n_1191));
   XNOR2_X1 i_1803 (.A(n_1194), .B(n_1193), .ZN(n_1192));
   NAND2_X1 i_1804 (.A1(A[19]), .A2(B[4]), .ZN(n_1193));
   NAND2_X1 i_1805 (.A1(A[20]), .A2(B[3]), .ZN(n_1194));
   INV_X1 i_1806 (.A(n_1197), .ZN(n_1196));
   XOR2_X1 i_1807 (.A(n_1212), .B(n_1198), .Z(n_1197));
   OAI22_X1 i_1808 (.A1(n_1209), .A2(n_1205), .B1(n_1200), .B2(n_1199), .ZN(
      n_1198));
   NAND2_X1 i_1809 (.A1(A[3]), .A2(B[20]), .ZN(n_1199));
   OAI21_X1 i_1810 (.A(n_1203), .B1(n_1209), .B2(n_1205), .ZN(n_1200));
   INV_X1 i_1811 (.A(n_1204), .ZN(n_1203));
   AOI22_X1 i_1812 (.A1(A[5]), .A2(B[18]), .B1(A[4]), .B2(B[19]), .ZN(n_1204));
   NAND2_X1 i_1813 (.A1(A[5]), .A2(B[19]), .ZN(n_1205));
   NAND2_X1 i_1814 (.A1(A[4]), .A2(B[18]), .ZN(n_1209));
   XNOR2_X1 i_1815 (.A(n_1222), .B(n_1213), .ZN(n_1212));
   AOI21_X1 i_1816 (.A(n_1221), .B1(n_1220), .B2(n_1214), .ZN(n_1213));
   NAND2_X1 i_1817 (.A1(A[9]), .A2(B[14]), .ZN(n_1214));
   OR3_X1 i_1818 (.A1(n_1235), .A2(n_229), .A3(n_1060), .ZN(n_1220));
   AOI22_X1 i_1819 (.A1(A[10]), .A2(B[13]), .B1(A[11]), .B2(B[12]), .ZN(n_1221));
   AOI21_X1 i_1820 (.A(n_1228), .B1(n_1226), .B2(n_1225), .ZN(n_1222));
   NOR2_X1 i_1821 (.A1(n_1232), .A2(n_170), .ZN(n_1225));
   NOR2_X1 i_1822 (.A1(n_1228), .A2(n_1227), .ZN(n_1226));
   AOI22_X1 i_1823 (.A1(A[8]), .A2(B[15]), .B1(A[7]), .B2(B[16]), .ZN(n_1227));
   NOR2_X1 i_1824 (.A1(n_1231), .A2(n_1230), .ZN(n_1228));
   NAND2_X1 i_1825 (.A1(A[8]), .A2(B[16]), .ZN(n_1230));
   NAND2_X1 i_1826 (.A1(A[7]), .A2(B[15]), .ZN(n_1231));
   INV_X1 i_1827 (.A(B[17]), .ZN(n_1232));
   INV_X1 i_1828 (.A(A[11]), .ZN(n_1235));
   XNOR2_X1 i_1829 (.A(n_1263), .B(n_1239), .ZN(n_1236));
   OAI22_X1 i_1830 (.A1(n_1262), .A2(n_1261), .B1(n_1260), .B2(n_1259), .ZN(
      n_1239));
   NAND2_X1 i_1831 (.A1(A[0]), .A2(B[23]), .ZN(n_1259));
   XNOR2_X1 i_1832 (.A(n_1262), .B(n_1261), .ZN(n_1260));
   NAND2_X1 i_1833 (.A1(A[1]), .A2(B[22]), .ZN(n_1261));
   NAND2_X1 i_1834 (.A1(A[2]), .A2(B[21]), .ZN(n_1262));
   AOI22_X1 i_1835 (.A1(n_1294), .A2(n_1293), .B1(n_1292), .B2(n_1266), .ZN(
      n_1263));
   INV_X1 i_1836 (.A(n_1266), .ZN(n_1264));
   OAI22_X1 i_1837 (.A1(n_1016), .A2(n_1157), .B1(n_1173), .B2(n_1290), .ZN(
      n_1266));
   NOR2_X1 i_1838 (.A1(n_1291), .A2(n_1290), .ZN(n_1289));
   AOI22_X1 i_1839 (.A1(A[13]), .A2(B[9]), .B1(A[14]), .B2(B[8]), .ZN(n_1290));
   NOR2_X1 i_1840 (.A1(n_1016), .A2(n_1157), .ZN(n_1291));
   XOR2_X1 i_1841 (.A(n_1294), .B(n_1293), .Z(n_1292));
   OAI21_X1 i_1842 (.A(n_1299), .B1(n_1296), .B2(n_1295), .ZN(n_1293));
   OAI21_X1 i_1843 (.A(n_1303), .B1(n_1301), .B2(n_1300), .ZN(n_1294));
   NAND2_X1 i_1844 (.A1(A[18]), .A2(B[4]), .ZN(n_1295));
   NAND2_X1 i_1845 (.A1(n_1299), .A2(n_1297), .ZN(n_1296));
   INV_X1 i_1846 (.A(n_1298), .ZN(n_1297));
   AOI22_X1 i_1847 (.A1(A[20]), .A2(B[2]), .B1(A[19]), .B2(B[3]), .ZN(n_1298));
   OR2_X1 i_1848 (.A1(n_954), .A2(n_1194), .ZN(n_1299));
   NAND2_X1 i_1849 (.A1(A[15]), .A2(B[7]), .ZN(n_1300));
   NAND2_X1 i_1850 (.A1(n_1303), .A2(n_1302), .ZN(n_1301));
   OAI22_X1 i_1851 (.A1(n_1305), .A2(n_169), .B1(n_1029), .B2(n_1027), .ZN(
      n_1302));
   OR3_X1 i_1852 (.A1(n_1152), .A2(n_1029), .A3(n_1305), .ZN(n_1303));
   INV_X1 i_1853 (.A(A[16]), .ZN(n_1305));
   INV_X1 i_1854 (.A(A[21]), .ZN(n_1317));
   NAND2_X1 i_1855 (.A1(B[4]), .A2(A[22]), .ZN(n_1318));
   NOR3_X1 i_1856 (.A1(n_1318), .A2(n_1317), .A3(n_424), .ZN(n_1319));
   AOI22_X1 i_1857 (.A1(B[3]), .A2(A[22]), .B1(B[4]), .B2(A[21]), .ZN(n_1320));
   NOR2_X1 i_1858 (.A1(n_1319), .A2(n_1320), .ZN(n_1321));
   INV_X1 i_1859 (.A(A[20]), .ZN(n_1322));
   NOR2_X1 i_1860 (.A1(n_1322), .A2(n_1029), .ZN(n_1323));
   XNOR2_X1 i_1861 (.A(n_1321), .B(n_1323), .ZN(n_1324));
   AOI22_X1 i_1862 (.A1(n_1190), .A2(n_1154), .B1(n_1153), .B2(n_1147), .ZN(
      n_1325));
   XNOR2_X1 i_1863 (.A(n_1324), .B(n_1325), .ZN(n_1326));
   AOI22_X1 i_1864 (.A1(A[21]), .A2(B[2]), .B1(B[0]), .B2(A[23]), .ZN(n_1327));
   NAND2_X1 i_1865 (.A1(B[2]), .A2(A[23]), .ZN(n_1328));
   NOR2_X1 i_1866 (.A1(n_1328), .A2(n_988), .ZN(n_1329));
   NOR2_X1 i_1867 (.A1(n_1328), .A2(n_949), .ZN(n_1330));
   INV_X1 i_1868 (.A(n_1329), .ZN(n_1331));
   AOI21_X1 i_1869 (.A(n_1327), .B1(n_1331), .B2(n_949), .ZN(n_1332));
   AOI22_X1 i_1870 (.A1(A[22]), .A2(B[2]), .B1(A[23]), .B2(B[1]), .ZN(n_1333));
   NOR2_X1 i_1871 (.A1(n_1330), .A2(n_1333), .ZN(n_1334));
   AOI21_X1 i_1872 (.A(n_1330), .B1(n_1332), .B2(n_1334), .ZN(n_1338));
   INV_X1 i_1873 (.A(A[10]), .ZN(n_1339));
   NAND2_X1 i_1874 (.A1(A[11]), .A2(B[14]), .ZN(n_1341));
   NAND2_X1 i_1875 (.A1(A[12]), .A2(B[12]), .ZN(n_1343));
   NAND2_X1 i_1876 (.A1(B[10]), .A2(A[15]), .ZN(n_1344));
   OR3_X1 i_1877 (.A1(n_1341), .A2(n_1339), .A3(n_229), .ZN(n_1345));
   OAI22_X1 i_1878 (.A1(n_1339), .A2(n_559), .B1(n_229), .B2(n_1235), .ZN(n_1346));
   NAND2_X1 i_1879 (.A1(n_1345), .A2(n_1346), .ZN(n_1348));
   OAI21_X1 i_1880 (.A(n_1345), .B1(n_1348), .B2(n_1343), .ZN(n_1349));
   NOR2_X1 i_1881 (.A1(n_1344), .A2(n_1157), .ZN(n_1357));
   INV_X1 i_1882 (.A(n_1357), .ZN(n_1358));
   AOI22_X1 i_1883 (.A1(A[14]), .A2(B[10]), .B1(A[15]), .B2(B[9]), .ZN(n_1359));
   OR2_X1 i_1884 (.A1(n_1357), .A2(n_1359), .ZN(n_1360));
   OAI21_X1 i_1885 (.A(n_1358), .B1(n_1360), .B2(n_1164), .ZN(n_1361));
   XOR2_X1 i_1886 (.A(n_1349), .B(n_1361), .Z(n_1362));
   NAND2_X1 i_1887 (.A1(A[9]), .A2(B[15]), .ZN(n_1363));
   XNOR2_X1 i_1888 (.A(n_1363), .B(n_1230), .ZN(n_1364));
   OAI33_X1 i_1889 (.A1(n_1364), .A2(n_556), .A3(n_1232), .B1(n_458), .B2(n_592), 
      .B3(n_1363), .ZN(n_1365));
   AOI22_X1 i_1890 (.A1(n_1365), .A2(n_1362), .B1(n_1361), .B2(n_1349), .ZN(
      n_1366));
   INV_X1 i_1891 (.A(B[21]), .ZN(n_1367));
   INV_X1 i_1892 (.A(B[22]), .ZN(n_1368));
   NAND4_X1 i_1893 (.A1(A[4]), .A2(A[3]), .A3(B[21]), .A4(B[22]), .ZN(n_1369));
   OAI22_X1 i_1894 (.A1(n_1367), .A2(n_422), .B1(n_1368), .B2(n_99), .ZN(n_1370));
   NAND2_X1 i_1895 (.A1(n_1369), .A2(n_1370), .ZN(n_1371));
   NAND2_X1 i_1896 (.A1(A[2]), .A2(B[23]), .ZN(n_1372));
   OAI21_X1 i_1897 (.A(n_1369), .B1(n_1371), .B2(n_1372), .ZN(n_1373));
   XNOR2_X1 i_1898 (.A(n_1366), .B(n_1373), .ZN(n_1374));
   NAND2_X1 i_1899 (.A1(B[7]), .A2(A[18]), .ZN(n_1375));
   NOR3_X1 i_1900 (.A1(n_1317), .A2(n_1194), .A3(n_340), .ZN(n_1376));
   INV_X1 i_1901 (.A(n_424), .ZN(n_1377));
   INV_X1 i_1902 (.A(n_340), .ZN(n_1378));
   AOI22_X1 i_1903 (.A1(n_1377), .A2(A[21]), .B1(n_1378), .B2(A[20]), .ZN(n_1381));
   NOR2_X1 i_1904 (.A1(n_1381), .A2(n_1376), .ZN(n_1382));
   AND2_X1 i_1905 (.A1(A[19]), .A2(B[5]), .ZN(n_1383));
   AOI21_X1 i_1906 (.A(n_1376), .B1(n_1382), .B2(n_1383), .ZN(n_1384));
   NOR2_X1 i_1907 (.A1(n_1375), .A2(n_1152), .ZN(n_1402));
   AOI22_X1 i_1908 (.A1(A[17]), .A2(B[7]), .B1(A[18]), .B2(B[6]), .ZN(n_1403));
   NOR2_X1 i_1909 (.A1(n_1402), .A2(n_1403), .ZN(n_1404));
   AND2_X1 i_1910 (.A1(A[16]), .A2(B[8]), .ZN(n_1405));
   AOI21_X1 i_1911 (.A(n_1402), .B1(n_1404), .B2(n_1405), .ZN(n_1406));
   XNOR2_X1 i_1912 (.A(n_1384), .B(n_1406), .ZN(n_1409));
   OAI22_X1 i_1913 (.A1(n_1409), .A2(n_1328), .B1(n_1384), .B2(n_1406), .ZN(
      n_1410));
   XOR2_X1 i_1914 (.A(n_1374), .B(n_1410), .Z(n_1411));
   OAI22_X1 i_1915 (.A1(n_1326), .A2(n_1338), .B1(n_1324), .B2(n_1325), .ZN(
      n_1412));
   XOR2_X1 i_1916 (.A(n_1411), .B(n_1412), .Z(n_1413));
   XOR2_X1 i_1917 (.A(n_1360), .B(n_1164), .Z(n_1414));
   XOR2_X1 i_1918 (.A(n_1348), .B(n_1343), .Z(n_1415));
   XOR2_X1 i_1919 (.A(n_1414), .B(n_1415), .Z(n_1418));
   NAND2_X1 i_1920 (.A1(A[7]), .A2(B[17]), .ZN(n_1419));
   XOR2_X1 i_1921 (.A(n_1364), .B(n_1419), .Z(n_1420));
   AOI22_X1 i_1922 (.A1(n_1418), .A2(n_1420), .B1(n_1414), .B2(n_1415), .ZN(
      n_1421));
   XNOR2_X1 i_1923 (.A(n_1409), .B(n_1328), .ZN(n_1422));
   XOR2_X1 i_1924 (.A(n_1421), .B(n_1422), .Z(n_1423));
   XOR2_X1 i_1925 (.A(n_1382), .B(n_1383), .Z(n_1424));
   XOR2_X1 i_1926 (.A(n_1404), .B(n_1405), .Z(n_1425));
   XOR2_X1 i_1927 (.A(n_1424), .B(n_1425), .Z(n_1426));
   XNOR2_X1 i_1928 (.A(n_1332), .B(n_1334), .ZN(n_1436));
   NAND2_X1 i_1929 (.A1(n_1426), .A2(n_1436), .ZN(n_1441));
   OAI21_X1 i_1930 (.A(n_1441), .B1(n_1425), .B2(n_1424), .ZN(n_1442));
   AOI22_X1 i_1931 (.A1(n_1423), .A2(n_1442), .B1(n_1421), .B2(n_1422), .ZN(
      n_1443));
   AOI22_X1 i_1932 (.A1(n_1413), .A2(n_1443), .B1(n_1411), .B2(n_1412), .ZN(
      n_1444));
   INV_X1 i_1933 (.A(n_1410), .ZN(n_1447));
   INV_X1 i_1934 (.A(n_1449), .ZN(n_1448));
   AOI22_X1 i_1935 (.A1(n_1453), .A2(n_1452), .B1(n_1502), .B2(n_1450), .ZN(
      n_1449));
   XOR2_X1 i_1936 (.A(n_1453), .B(n_1452), .Z(n_1450));
   XOR2_X1 i_1937 (.A(n_1455), .B(n_1454), .Z(n_1452));
   OAI22_X1 i_1938 (.A1(n_1477), .A2(n_1476), .B1(n_1501), .B2(n_1461), .ZN(
      n_1453));
   NOR2_X1 i_1939 (.A1(n_1533), .A2(n_99), .ZN(n_1454));
   NOR2_X1 i_1940 (.A1(n_1459), .A2(n_1456), .ZN(n_1455));
   AOI22_X1 i_1941 (.A1(A[5]), .A2(B[21]), .B1(A[4]), .B2(B[22]), .ZN(n_1456));
   NOR3_X1 i_1942 (.A1(n_422), .A2(n_1460), .A3(n_1367), .ZN(n_1459));
   NAND2_X1 i_1943 (.A1(A[5]), .A2(B[22]), .ZN(n_1460));
   XNOR2_X1 i_1944 (.A(n_1477), .B(n_1476), .ZN(n_1461));
   OAI21_X1 i_1945 (.A(n_1481), .B1(n_1480), .B2(n_1478), .ZN(n_1476));
   OAI21_X1 i_1946 (.A(n_1485), .B1(n_1483), .B2(n_1482), .ZN(n_1477));
   NOR2_X1 i_1947 (.A1(n_422), .A2(n_856), .ZN(n_1478));
   INV_X1 i_1948 (.A(n_1480), .ZN(n_1479));
   NOR3_X1 i_1949 (.A1(n_1205), .A2(n_170), .A3(n_1532), .ZN(n_1480));
   OAI21_X1 i_1950 (.A(n_1205), .B1(n_1532), .B2(n_170), .ZN(n_1481));
   NOR2_X1 i_1951 (.A1(n_1534), .A2(n_1533), .ZN(n_1482));
   INV_X1 i_1952 (.A(n_1484), .ZN(n_1483));
   NAND3_X1 i_1953 (.A1(A[3]), .A2(n_1530), .A3(B[22]), .ZN(n_1484));
   OAI22_X1 i_1954 (.A1(n_99), .A2(n_1367), .B1(n_33), .B2(n_1368), .ZN(n_1485));
   AOI22_X1 i_1955 (.A1(n_1212), .A2(n_1198), .B1(n_1531), .B2(n_1213), .ZN(
      n_1501));
   XOR2_X1 i_1956 (.A(n_1509), .B(n_1503), .Z(n_1502));
   OAI22_X1 i_1957 (.A1(n_1205), .A2(n_1508), .B1(n_1505), .B2(n_1504), .ZN(
      n_1503));
   NAND2_X1 i_1958 (.A1(A[7]), .A2(B[18]), .ZN(n_1504));
   OAI21_X1 i_1959 (.A(n_1506), .B1(n_1205), .B2(n_1508), .ZN(n_1505));
   INV_X1 i_1960 (.A(n_1507), .ZN(n_1506));
   AOI22_X1 i_1961 (.A1(A[5]), .A2(B[20]), .B1(A[6]), .B2(B[19]), .ZN(n_1507));
   NAND2_X1 i_1962 (.A1(A[6]), .A2(B[20]), .ZN(n_1508));
   XOR2_X1 i_1963 (.A(n_1525), .B(n_1521), .Z(n_1509));
   OAI33_X1 i_1964 (.A1(n_458), .A2(n_1232), .A3(n_1522), .B1(n_1363), .B2(
      n_1339), .B3(n_592), .ZN(n_1521));
   XNOR2_X1 i_1965 (.A(n_1524), .B(n_1523), .ZN(n_1522));
   NAND2_X1 i_1966 (.A1(A[10]), .A2(B[15]), .ZN(n_1523));
   NAND2_X1 i_1967 (.A1(A[9]), .A2(B[16]), .ZN(n_1524));
   OAI22_X1 i_1968 (.A1(n_1343), .A2(n_1529), .B1(n_1341), .B2(n_1526), .ZN(
      n_1525));
   OAI21_X1 i_1969 (.A(n_1527), .B1(n_1343), .B2(n_1529), .ZN(n_1526));
   INV_X1 i_1970 (.A(n_1528), .ZN(n_1527));
   AOI22_X1 i_1971 (.A1(A[13]), .A2(B[12]), .B1(A[12]), .B2(B[13]), .ZN(n_1528));
   NAND2_X1 i_1972 (.A1(A[13]), .A2(B[13]), .ZN(n_1529));
   INV_X1 i_1973 (.A(n_1262), .ZN(n_1530));
   INV_X1 i_1974 (.A(n_1222), .ZN(n_1531));
   INV_X1 i_1975 (.A(B[18]), .ZN(n_1532));
   INV_X1 i_1976 (.A(B[23]), .ZN(n_1533));
   INV_X1 i_1977 (.A(A[1]), .ZN(n_1534));
   XNOR2_X1 i_1978 (.A(n_1574), .B(n_1553), .ZN(n_1535));
   XOR2_X1 i_1979 (.A(n_1563), .B(n_1554), .Z(n_1553));
   XOR2_X1 i_1980 (.A(n_1557), .B(n_1555), .Z(n_1554));
   NAND2_X1 i_1981 (.A1(n_1560), .A2(n_1558), .ZN(n_1555));
   NAND2_X1 i_1982 (.A1(B[20]), .A2(A[9]), .ZN(n_1557));
   OR2_X1 i_1983 (.A1(n_1562), .A2(n_1561), .ZN(n_1558));
   INV_X1 i_1984 (.A(n_1560), .ZN(n_1559));
   NAND2_X1 i_1985 (.A1(n_1562), .A2(n_1561), .ZN(n_1560));
   NAND2_X1 i_1986 (.A1(B[19]), .A2(A[10]), .ZN(n_1561));
   NAND2_X1 i_1987 (.A1(B[18]), .A2(A[11]), .ZN(n_1562));
   XOR2_X1 i_1988 (.A(n_1567), .B(n_1566), .Z(n_1563));
   NAND2_X1 i_1989 (.A1(n_1569), .A2(n_1568), .ZN(n_1566));
   NAND2_X1 i_1990 (.A1(B[23]), .A2(A[6]), .ZN(n_1567));
   OAI22_X1 i_1991 (.A1(n_1367), .A2(n_458), .B1(n_556), .B2(n_1368), .ZN(n_1568));
   NAND3_X1 i_1992 (.A1(A[8]), .A2(n_1573), .A3(B[22]), .ZN(n_1569));
   NOR2_X1 i_1993 (.A1(n_1367), .A2(n_556), .ZN(n_1573));
   AOI22_X1 i_1994 (.A1(n_1610), .A2(n_1609), .B1(n_1608), .B2(n_1575), .ZN(
      n_1574));
   AOI22_X1 i_1995 (.A1(n_1586), .A2(n_1580), .B1(n_1579), .B2(n_1576), .ZN(
      n_1575));
   INV_X1 i_1996 (.A(n_1577), .ZN(n_1576));
   AOI21_X1 i_1997 (.A(n_1459), .B1(n_1455), .B2(n_1454), .ZN(n_1577));
   XOR2_X1 i_1998 (.A(n_1586), .B(n_1580), .Z(n_1579));
   OAI22_X1 i_1999 (.A1(n_1504), .A2(n_1590), .B1(n_1508), .B2(n_1588), .ZN(
      n_1580));
   OAI21_X1 i_2000 (.A(n_1601), .B1(n_1524), .B2(n_1607), .ZN(n_1586));
   NOR2_X1 i_2001 (.A1(n_1589), .A2(n_1588), .ZN(n_1587));
   AOI22_X1 i_2002 (.A1(B[19]), .A2(A[7]), .B1(B[18]), .B2(A[8]), .ZN(n_1588));
   NOR2_X1 i_2003 (.A1(n_1504), .A2(n_1590), .ZN(n_1589));
   NAND2_X1 i_2004 (.A1(B[19]), .A2(A[8]), .ZN(n_1590));
   NAND2_X1 i_2005 (.A1(n_1604), .A2(n_1602), .ZN(n_1601));
   INV_X1 i_2006 (.A(n_1603), .ZN(n_1602));
   NAND2_X1 i_2007 (.A1(B[15]), .A2(A[11]), .ZN(n_1603));
   NOR2_X1 i_2008 (.A1(n_1606), .A2(n_1605), .ZN(n_1604));
   AOI22_X1 i_2009 (.A1(B[17]), .A2(A[9]), .B1(B[16]), .B2(A[10]), .ZN(n_1605));
   NOR2_X1 i_2010 (.A1(n_1524), .A2(n_1607), .ZN(n_1606));
   NAND2_X1 i_2011 (.A1(B[17]), .A2(A[10]), .ZN(n_1607));
   XOR2_X1 i_2012 (.A(n_1610), .B(n_1609), .Z(n_1608));
   AOI22_X1 i_2013 (.A1(n_1649), .A2(n_1613), .B1(n_1612), .B2(n_1611), .ZN(
      n_1609));
   AOI21_X1 i_2014 (.A(n_1622), .B1(n_1621), .B2(n_1614), .ZN(n_1610));
   NOR2_X1 i_2015 (.A1(n_422), .A2(n_1533), .ZN(n_1611));
   XOR2_X1 i_2016 (.A(n_1649), .B(n_1613), .Z(n_1612));
   NOR2_X1 i_2017 (.A1(n_170), .A2(n_1367), .ZN(n_1613));
   OAI22_X1 i_2018 (.A1(n_1529), .A2(n_1617), .B1(n_1616), .B2(n_1615), .ZN(
      n_1614));
   NAND2_X1 i_2019 (.A1(B[14]), .A2(A[12]), .ZN(n_1615));
   XNOR2_X1 i_2020 (.A(n_1529), .B(n_1617), .ZN(n_1616));
   NAND2_X1 i_2021 (.A1(B[12]), .A2(A[14]), .ZN(n_1617));
   INV_X1 i_2022 (.A(n_1621), .ZN(n_1620));
   AOI21_X1 i_2023 (.A(n_1622), .B1(n_1624), .B2(n_1623), .ZN(n_1621));
   NOR2_X1 i_2024 (.A1(n_1624), .A2(n_1623), .ZN(n_1622));
   AOI21_X1 i_2025 (.A(n_1629), .B1(n_1627), .B2(n_1626), .ZN(n_1623));
   AOI21_X1 i_2026 (.A(n_1647), .B1(n_1636), .B2(n_1634), .ZN(n_1624));
   AND2_X1 i_2027 (.A1(B[11]), .A2(A[15]), .ZN(n_1626));
   NOR2_X1 i_2028 (.A1(n_1629), .A2(n_1628), .ZN(n_1627));
   AOI22_X1 i_2029 (.A1(B[10]), .A2(A[16]), .B1(B[9]), .B2(A[17]), .ZN(n_1628));
   NOR2_X1 i_2030 (.A1(n_1631), .A2(n_1630), .ZN(n_1629));
   NAND2_X1 i_2031 (.A1(B[10]), .A2(A[17]), .ZN(n_1630));
   NAND2_X1 i_2032 (.A1(B[9]), .A2(A[16]), .ZN(n_1631));
   INV_X1 i_2033 (.A(n_1635), .ZN(n_1634));
   NAND2_X1 i_2034 (.A1(B[6]), .A2(A[20]), .ZN(n_1635));
   NOR2_X1 i_2035 (.A1(n_1647), .A2(n_1640), .ZN(n_1636));
   AOI22_X1 i_2036 (.A1(B[8]), .A2(A[18]), .B1(B[7]), .B2(A[19]), .ZN(n_1640));
   NOR2_X1 i_2037 (.A1(n_1375), .A2(n_1648), .ZN(n_1647));
   NAND2_X1 i_2038 (.A1(B[8]), .A2(A[19]), .ZN(n_1648));
   INV_X1 i_2039 (.A(n_1460), .ZN(n_1649));
   XNOR2_X1 i_2040 (.A(n_1579), .B(n_1577), .ZN(n_1650));
   INV_X1 i_2041 (.A(n_1373), .ZN(n_1652));
   INV_X1 i_2042 (.A(n_1374), .ZN(n_1653));
   OAI22_X1 i_2043 (.A1(n_1652), .A2(n_1366), .B1(n_1653), .B2(n_1447), .ZN(
      n_1654));
   XOR2_X1 i_2044 (.A(n_1650), .B(n_1654), .Z(n_1655));
   XNOR2_X1 i_2045 (.A(n_1620), .B(n_1614), .ZN(n_1658));
   AOI22_X1 i_2046 (.A1(n_1655), .A2(n_1658), .B1(n_1650), .B2(n_1654), .ZN(
      n_1659));
   XOR2_X1 i_2047 (.A(n_1608), .B(n_1575), .Z(n_1660));
   NOR2_X1 i_2048 (.A1(n_1659), .A2(n_1660), .ZN(n_1661));
   AOI21_X1 i_2049 (.A(n_1661), .B1(n_1659), .B2(n_1660), .ZN(n_1662));
   INV_X1 i_2050 (.A(B[12]), .ZN(n_1676));
   NAND2_X1 i_2051 (.A1(B[13]), .A2(A[16]), .ZN(n_1698));
   OR3_X1 i_2052 (.A1(n_1698), .A2(n_1676), .A3(n_558), .ZN(n_1699));
   OAI22_X1 i_2053 (.A1(n_1676), .A2(n_1305), .B1(n_558), .B2(n_229), .ZN(n_1700));
   NAND2_X1 i_2054 (.A1(n_1699), .A2(n_1700), .ZN(n_1701));
   NAND2_X1 i_2055 (.A1(B[14]), .A2(A[14]), .ZN(n_1702));
   XNOR2_X1 i_2056 (.A(n_1701), .B(n_1702), .ZN(n_1703));
   NAND2_X1 i_2057 (.A1(B[16]), .A2(A[12]), .ZN(n_1704));
   NAND2_X1 i_2058 (.A1(B[17]), .A2(A[11]), .ZN(n_1705));
   XNOR2_X1 i_2059 (.A(n_1704), .B(n_1705), .ZN(n_1706));
   NAND2_X1 i_2060 (.A1(B[15]), .A2(A[13]), .ZN(n_1707));
   XNOR2_X1 i_2061 (.A(n_1706), .B(n_1707), .ZN(n_1708));
   XOR2_X1 i_2062 (.A(n_1708), .B(n_1703), .Z(n_1709));
   NAND2_X1 i_2063 (.A1(A[9]), .A2(B[18]), .ZN(n_1710));
   INV_X1 i_2064 (.A(B[19]), .ZN(n_1711));
   NOR3_X1 i_2065 (.A1(n_1710), .A2(n_1711), .A3(n_1339), .ZN(n_1712));
   AOI22_X1 i_2066 (.A1(B[19]), .A2(A[9]), .B1(B[18]), .B2(A[10]), .ZN(n_1713));
   NOR2_X1 i_2067 (.A1(n_1712), .A2(n_1713), .ZN(n_1714));
   NOR2_X1 i_2068 (.A1(n_458), .A2(n_856), .ZN(n_1715));
   XNOR2_X1 i_2069 (.A(n_1714), .B(n_1715), .ZN(n_1716));
   XNOR2_X1 i_2070 (.A(n_1709), .B(n_1716), .ZN(n_1717));
   AOI21_X1 i_2071 (.A(n_1661), .B1(n_1717), .B2(n_1662), .ZN(n_1718));
   XOR2_X1 i_2072 (.A(n_1757), .B(n_1720), .Z(n_1719));
   XOR2_X1 i_2073 (.A(n_1728), .B(n_1721), .Z(n_1720));
   XNOR2_X1 i_2074 (.A(n_1723), .B(n_1722), .ZN(n_1721));
   NOR2_X1 i_2075 (.A1(n_1792), .A2(n_169), .ZN(n_1722));
   NOR2_X1 i_2076 (.A1(n_1725), .A2(n_1724), .ZN(n_1723));
   AOI22_X1 i_2077 (.A1(B[7]), .A2(A[22]), .B1(B[8]), .B2(A[21]), .ZN(n_1724));
   NOR2_X1 i_2078 (.A1(n_1783), .A2(n_1726), .ZN(n_1725));
   NAND2_X1 i_2079 (.A1(B[8]), .A2(A[22]), .ZN(n_1726));
   AOI22_X1 i_2080 (.A1(n_1737), .A2(n_1736), .B1(n_1734), .B2(n_1730), .ZN(
      n_1728));
   OAI21_X1 i_2081 (.A(n_1732), .B1(n_1710), .B2(n_1731), .ZN(n_1730));
   OAI21_X1 i_2082 (.A(n_1732), .B1(n_1790), .B2(n_1733), .ZN(n_1731));
   NAND2_X1 i_2083 (.A1(n_1790), .A2(n_1733), .ZN(n_1732));
   NOR2_X1 i_2084 (.A1(n_556), .A2(n_856), .ZN(n_1733));
   XOR2_X1 i_2085 (.A(n_1737), .B(n_1736), .Z(n_1734));
   OAI21_X1 i_2086 (.A(n_1740), .B1(n_1739), .B2(n_1738), .ZN(n_1736));
   OAI21_X1 i_2087 (.A(n_1745), .B1(n_1603), .B2(n_1704), .ZN(n_1737));
   NAND2_X1 i_2088 (.A1(B[14]), .A2(A[13]), .ZN(n_1738));
   OAI21_X1 i_2089 (.A(n_1740), .B1(n_1744), .B2(n_1743), .ZN(n_1739));
   NAND2_X1 i_2090 (.A1(n_1744), .A2(n_1743), .ZN(n_1740));
   NOR2_X1 i_2091 (.A1(n_229), .A2(n_557), .ZN(n_1743));
   NOR2_X1 i_2092 (.A1(n_1676), .A2(n_558), .ZN(n_1744));
   NAND2_X1 i_2093 (.A1(n_1791), .A2(n_1746), .ZN(n_1745));
   NOR2_X1 i_2094 (.A1(n_1755), .A2(n_1754), .ZN(n_1746));
   AOI22_X1 i_2095 (.A1(B[15]), .A2(A[12]), .B1(B[16]), .B2(A[11]), .ZN(n_1754));
   NOR2_X1 i_2096 (.A1(n_1603), .A2(n_1704), .ZN(n_1755));
   AOI22_X1 i_2097 (.A1(n_1786), .A2(n_1785), .B1(n_1784), .B2(n_1761), .ZN(
      n_1757));
   INV_X1 i_2098 (.A(n_1761), .ZN(n_1760));
   OAI22_X1 i_2099 (.A1(n_1635), .A2(n_1783), .B1(n_1648), .B2(n_1763), .ZN(
      n_1761));
   NOR2_X1 i_2100 (.A1(n_1782), .A2(n_1763), .ZN(n_1762));
   AOI22_X1 i_2101 (.A1(B[6]), .A2(A[21]), .B1(B[7]), .B2(A[20]), .ZN(n_1763));
   NOR2_X1 i_2102 (.A1(n_1635), .A2(n_1783), .ZN(n_1782));
   NAND2_X1 i_2103 (.A1(B[7]), .A2(A[21]), .ZN(n_1783));
   XOR2_X1 i_2104 (.A(n_1786), .B(n_1785), .Z(n_1784));
   OAI22_X1 i_2105 (.A1(n_1630), .A2(n_1789), .B1(n_1788), .B2(n_1787), .ZN(
      n_1785));
   NOR2_X1 i_2106 (.A1(n_1792), .A2(n_1029), .ZN(n_1786));
   NAND2_X1 i_2107 (.A1(B[9]), .A2(A[18]), .ZN(n_1787));
   XNOR2_X1 i_2108 (.A(n_1630), .B(n_1789), .ZN(n_1788));
   NAND2_X1 i_2109 (.A1(B[11]), .A2(A[16]), .ZN(n_1789));
   INV_X1 i_2110 (.A(n_1590), .ZN(n_1790));
   INV_X1 i_2111 (.A(n_1607), .ZN(n_1791));
   INV_X1 i_2112 (.A(A[23]), .ZN(n_1792));
   XOR2_X1 i_2113 (.A(n_1812), .B(n_1794), .Z(n_1793));
   XNOR2_X1 i_2114 (.A(n_1796), .B(n_1795), .ZN(n_1794));
   AOI22_X1 i_2115 (.A1(n_1574), .A2(n_1553), .B1(n_1563), .B2(n_1554), .ZN(
      n_1795));
   XOR2_X1 i_2116 (.A(n_1811), .B(n_1797), .Z(n_1796));
   AOI21_X1 i_2117 (.A(n_1807), .B1(n_1806), .B2(n_1805), .ZN(n_1797));
   XNOR2_X1 i_2118 (.A(n_1845), .B(n_1844), .ZN(n_1805));
   AOI21_X1 i_2119 (.A(n_1807), .B1(n_1810), .B2(n_1808), .ZN(n_1806));
   NOR2_X1 i_2120 (.A1(n_1810), .A2(n_1808), .ZN(n_1807));
   XOR2_X1 i_2121 (.A(n_1851), .B(n_1809), .Z(n_1808));
   NAND2_X1 i_2122 (.A1(B[14]), .A2(A[15]), .ZN(n_1809));
   XOR2_X1 i_2123 (.A(n_1869), .B(n_1868), .Z(n_1810));
   AOI22_X1 i_2124 (.A1(n_1720), .A2(n_1757), .B1(n_1728), .B2(n_1721), .ZN(
      n_1811));
   XOR2_X1 i_2125 (.A(n_1832), .B(n_1813), .Z(n_1812));
   XOR2_X1 i_2126 (.A(n_1823), .B(n_1814), .Z(n_1813));
   XOR2_X1 i_2127 (.A(n_1822), .B(n_1815), .Z(n_1814));
   AOI21_X1 i_2128 (.A(n_1559), .B1(n_1558), .B2(n_1557), .ZN(n_1815));
   INV_X1 i_2129 (.A(n_1822), .ZN(n_1821));
   AOI21_X1 i_2130 (.A(n_1875), .B1(n_1567), .B2(n_1569), .ZN(n_1822));
   OAI22_X1 i_2131 (.A1(n_1830), .A2(n_1829), .B1(n_1828), .B2(n_1824), .ZN(
      n_1823));
   AOI21_X1 i_2132 (.A(n_1827), .B1(n_1573), .B2(n_1825), .ZN(n_1824));
   NOR2_X1 i_2133 (.A1(n_1827), .A2(n_1826), .ZN(n_1825));
   AOI22_X1 i_2134 (.A1(B[23]), .A2(A[5]), .B1(B[22]), .B2(A[6]), .ZN(n_1826));
   NOR2_X1 i_2135 (.A1(n_1460), .A2(n_1567), .ZN(n_1827));
   XNOR2_X1 i_2136 (.A(n_1830), .B(n_1829), .ZN(n_1828));
   AOI21_X1 i_2137 (.A(n_1712), .B1(n_1714), .B2(n_1715), .ZN(n_1829));
   INV_X1 i_2138 (.A(n_1831), .ZN(n_1830));
   OAI22_X1 i_2139 (.A1(n_1707), .A2(n_1706), .B1(n_1704), .B2(n_1705), .ZN(
      n_1831));
   XOR2_X1 i_2140 (.A(n_1842), .B(n_1833), .Z(n_1832));
   XNOR2_X1 i_2141 (.A(n_1841), .B(n_1834), .ZN(n_1833));
   NOR2_X1 i_2142 (.A1(n_1839), .A2(n_1837), .ZN(n_1834));
   AOI22_X1 i_2143 (.A1(B[21]), .A2(A[9]), .B1(B[22]), .B2(A[8]), .ZN(n_1837));
   INV_X1 i_2144 (.A(n_1839), .ZN(n_1838));
   NOR3_X1 i_2145 (.A1(n_458), .A2(n_1840), .A3(n_1367), .ZN(n_1839));
   NAND2_X1 i_2146 (.A1(B[22]), .A2(A[9]), .ZN(n_1840));
   NAND2_X1 i_2147 (.A1(B[23]), .A2(A[7]), .ZN(n_1841));
   XOR2_X1 i_2148 (.A(n_1849), .B(n_1843), .Z(n_1842));
   OAI22_X1 i_2149 (.A1(n_1707), .A2(n_1848), .B1(n_1845), .B2(n_1844), .ZN(
      n_1843));
   NAND2_X1 i_2150 (.A1(B[17]), .A2(A[12]), .ZN(n_1844));
   OAI21_X1 i_2151 (.A(n_1846), .B1(n_1707), .B2(n_1848), .ZN(n_1845));
   INV_X1 i_2152 (.A(n_1847), .ZN(n_1846));
   AOI22_X1 i_2153 (.A1(B[16]), .A2(A[13]), .B1(B[15]), .B2(A[14]), .ZN(n_1847));
   NAND2_X1 i_2154 (.A1(B[16]), .A2(A[14]), .ZN(n_1848));
   XOR2_X1 i_2155 (.A(n_1853), .B(n_1850), .Z(n_1849));
   OAI33_X1 i_2156 (.A1(n_559), .A2(n_558), .A3(n_1851), .B1(n_229), .B2(n_1305), 
      .B3(n_1852), .ZN(n_1850));
   XNOR2_X1 i_2157 (.A(n_1698), .B(n_1852), .ZN(n_1851));
   NAND2_X1 i_2158 (.A1(B[12]), .A2(A[17]), .ZN(n_1852));
   OAI21_X1 i_2159 (.A(n_1870), .B1(n_1869), .B2(n_1868), .ZN(n_1853));
   NAND2_X1 i_2160 (.A1(B[11]), .A2(A[18]), .ZN(n_1868));
   OAI21_X1 i_2161 (.A(n_1870), .B1(n_1872), .B2(n_1871), .ZN(n_1869));
   NAND2_X1 i_2162 (.A1(n_1872), .A2(n_1871), .ZN(n_1870));
   AND2_X1 i_2163 (.A1(B[10]), .A2(A[19]), .ZN(n_1871));
   AND2_X1 i_2164 (.A1(B[9]), .A2(A[20]), .ZN(n_1872));
   NAND2_X1 i_2165 (.A1(B[10]), .A2(A[20]), .ZN(n_1873));
   NAND2_X1 i_2166 (.A1(B[9]), .A2(A[19]), .ZN(n_1874));
   INV_X1 i_2167 (.A(n_1568), .ZN(n_1875));
   NAND2_X1 i_2168 (.A1(B[10]), .A2(A[18]), .ZN(n_1876));
   XNOR2_X1 i_2169 (.A(n_1876), .B(n_1874), .ZN(n_1877));
   NAND2_X1 i_2170 (.A1(B[11]), .A2(A[17]), .ZN(n_1878));
   OAI22_X1 i_2171 (.A1(n_1877), .A2(n_1878), .B1(n_1876), .B2(n_1874), .ZN(
      n_1879));
   OAI21_X1 i_2172 (.A(n_1783), .B1(n_425), .B2(n_1322), .ZN(n_1880));
   INV_X1 i_2173 (.A(A[22]), .ZN(n_1881));
   NOR2_X1 i_2174 (.A1(n_1881), .A2(n_169), .ZN(n_1882));
   NOR3_X1 i_2175 (.A1(n_1783), .A2(n_425), .A3(n_1322), .ZN(n_1883));
   OAI21_X1 i_2176 (.A(n_1880), .B1(n_1883), .B2(n_1882), .ZN(n_1884));
   OAI21_X1 i_2177 (.A(n_1699), .B1(n_1701), .B2(n_1702), .ZN(n_1885));
   XNOR2_X1 i_2178 (.A(n_1879), .B(n_1884), .ZN(n_1886));
   XNOR2_X1 i_2179 (.A(n_1886), .B(n_1885), .ZN(n_1887));
   XNOR2_X1 i_2180 (.A(n_1828), .B(n_1824), .ZN(n_1888));
   XOR2_X1 i_2181 (.A(n_1887), .B(n_1888), .Z(n_1889));
   AOI22_X1 i_2182 (.A1(n_1709), .A2(n_1716), .B1(n_1703), .B2(n_1708), .ZN(
      n_1890));
   NAND2_X1 i_2183 (.A1(n_1889), .A2(n_1890), .ZN(n_1891));
   OAI21_X1 i_2184 (.A(n_1891), .B1(n_1888), .B2(n_1887), .ZN(n_1892));
   INV_X1 i_2185 (.A(n_1883), .ZN(n_1893));
   AOI21_X1 i_2186 (.A(n_1896), .B1(n_1930), .B2(n_1895), .ZN(n_1894));
   AOI21_X1 i_2187 (.A(n_1896), .B1(n_1905), .B2(n_1897), .ZN(n_1895));
   NOR2_X1 i_2188 (.A1(n_1905), .A2(n_1897), .ZN(n_1896));
   XOR2_X1 i_2189 (.A(n_1907), .B(n_1906), .Z(n_1897));
   AOI21_X1 i_2190 (.A(n_1915), .B1(n_1914), .B2(n_1910), .ZN(n_1905));
   OAI22_X1 i_2191 (.A1(n_1873), .A2(n_1954), .B1(n_1951), .B2(n_1941), .ZN(
      n_1906));
   XNOR2_X1 i_2192 (.A(n_1909), .B(n_1908), .ZN(n_1907));
   NOR2_X1 i_2193 (.A1(n_1792), .A2(n_425), .ZN(n_1908));
   NOR2_X1 i_2194 (.A1(n_1923), .A2(n_1918), .ZN(n_1909));
   XNOR2_X1 i_2195 (.A(n_1912), .B(n_1911), .ZN(n_1910));
   NAND2_X1 i_2196 (.A1(B[15]), .A2(A[15]), .ZN(n_1911));
   XNOR2_X1 i_2197 (.A(n_1848), .B(n_1913), .ZN(n_1912));
   NAND2_X1 i_2198 (.A1(B[17]), .A2(A[13]), .ZN(n_1913));
   AOI21_X1 i_2199 (.A(n_1915), .B1(n_1917), .B2(n_1916), .ZN(n_1914));
   NOR2_X1 i_2200 (.A1(n_1917), .A2(n_1916), .ZN(n_1915));
   XOR2_X1 i_2201 (.A(n_1926), .B(n_1925), .Z(n_1916));
   AOI21_X1 i_2202 (.A(n_1918), .B1(n_1921), .B2(n_1920), .ZN(n_1917));
   NOR2_X1 i_2203 (.A1(n_1921), .A2(n_1920), .ZN(n_1918));
   OR2_X1 i_2204 (.A1(n_559), .A2(n_1305), .ZN(n_1920));
   OR2_X1 i_2205 (.A1(n_1923), .A2(n_1922), .ZN(n_1921));
   AOI22_X1 i_2206 (.A1(B[13]), .A2(A[17]), .B1(B[12]), .B2(A[18]), .ZN(n_1922));
   NOR2_X1 i_2207 (.A1(n_1852), .A2(n_1924), .ZN(n_1923));
   NAND2_X1 i_2208 (.A1(B[13]), .A2(A[18]), .ZN(n_1924));
   NOR2_X1 i_2209 (.A1(n_1339), .A2(n_856), .ZN(n_1925));
   NOR2_X1 i_2210 (.A1(n_1928), .A2(n_1927), .ZN(n_1926));
   AOI22_X1 i_2211 (.A1(B[19]), .A2(A[11]), .B1(B[18]), .B2(A[12]), .ZN(n_1927));
   NOR3_X1 i_2212 (.A1(n_1235), .A2(n_1929), .A3(n_1532), .ZN(n_1928));
   NAND2_X1 i_2213 (.A1(B[19]), .A2(A[12]), .ZN(n_1929));
   AOI22_X1 i_2214 (.A1(n_1952), .A2(n_1936), .B1(n_1935), .B2(n_1931), .ZN(
      n_1930));
   XNOR2_X1 i_2215 (.A(n_1726), .B(n_1932), .ZN(n_1931));
   XNOR2_X1 i_2216 (.A(n_1934), .B(n_1933), .ZN(n_1932));
   NOR2_X1 i_2217 (.A1(n_1955), .A2(n_1792), .ZN(n_1933));
   AOI21_X1 i_2218 (.A(n_1725), .B1(n_1723), .B2(n_1722), .ZN(n_1934));
   XOR2_X1 i_2219 (.A(n_1952), .B(n_1936), .Z(n_1935));
   XOR2_X1 i_2220 (.A(n_1951), .B(n_1941), .Z(n_1936));
   NAND2_X1 i_2221 (.A1(B[11]), .A2(A[19]), .ZN(n_1941));
   XNOR2_X1 i_2222 (.A(n_1873), .B(n_1954), .ZN(n_1951));
   OAI21_X1 i_2223 (.A(n_1953), .B1(n_1884), .B2(n_1956), .ZN(n_1952));
   NAND2_X1 i_2224 (.A1(n_1886), .A2(n_1885), .ZN(n_1953));
   NAND2_X1 i_2225 (.A1(B[9]), .A2(A[21]), .ZN(n_1954));
   INV_X1 i_2226 (.A(B[7]), .ZN(n_1955));
   INV_X1 i_2227 (.A(n_1879), .ZN(n_1956));
   NAND2_X1 i_2228 (.A1(B[18]), .A2(A[14]), .ZN(n_1957));
   NAND2_X1 i_2229 (.A1(A[13]), .A2(B[20]), .ZN(n_1958));
   NOR2_X1 i_2230 (.A1(n_1958), .A2(n_1929), .ZN(n_1959));
   AOI22_X1 i_2231 (.A1(B[19]), .A2(A[13]), .B1(B[20]), .B2(A[12]), .ZN(n_1960));
   NOR2_X1 i_2232 (.A1(n_1959), .A2(n_1960), .ZN(n_1961));
   XOR2_X1 i_2233 (.A(n_1961), .B(n_1957), .Z(n_1962));
   NAND2_X1 i_2234 (.A1(B[17]), .A2(A[15]), .ZN(n_1963));
   NAND2_X1 i_2235 (.A1(B[15]), .A2(A[16]), .ZN(n_1964));
   NAND2_X1 i_2236 (.A1(A[17]), .A2(B[16]), .ZN(n_1965));
   NOR2_X1 i_2237 (.A1(n_1964), .A2(n_1965), .ZN(n_1966));
   AOI22_X1 i_2238 (.A1(B[15]), .A2(A[17]), .B1(B[16]), .B2(A[16]), .ZN(n_1967));
   NOR2_X1 i_2239 (.A1(n_1966), .A2(n_1967), .ZN(n_1974));
   XOR2_X1 i_2240 (.A(n_1974), .B(n_1963), .Z(n_1975));
   XOR2_X1 i_2241 (.A(n_1962), .B(n_1975), .Z(n_1976));
   NAND2_X1 i_2242 (.A1(B[21]), .A2(A[11]), .ZN(n_1977));
   NAND2_X1 i_2243 (.A1(B[22]), .A2(A[10]), .ZN(n_1978));
   XNOR2_X1 i_2244 (.A(n_1977), .B(n_1978), .ZN(n_1979));
   NAND2_X1 i_2245 (.A1(B[23]), .A2(A[9]), .ZN(n_1980));
   XNOR2_X1 i_2246 (.A(n_1979), .B(n_1980), .ZN(n_1981));
   INV_X1 i_2247 (.A(n_1909), .ZN(n_1982));
   AOI22_X1 i_2248 (.A1(n_1982), .A2(n_1908), .B1(n_1907), .B2(n_1906), .ZN(
      n_1984));
   NAND2_X1 i_2249 (.A1(B[12]), .A2(A[20]), .ZN(n_1985));
   NAND2_X1 i_2250 (.A1(B[13]), .A2(A[19]), .ZN(n_1986));
   XNOR2_X1 i_2251 (.A(n_1985), .B(n_1986), .ZN(n_1987));
   NAND2_X1 i_2252 (.A1(B[14]), .A2(A[18]), .ZN(n_1988));
   XOR2_X1 i_2253 (.A(n_1987), .B(n_1988), .Z(n_1990));
   XNOR2_X1 i_2254 (.A(n_1990), .B(n_1984), .ZN(n_1991));
   NAND2_X1 i_2255 (.A1(B[10]), .A2(A[22]), .ZN(n_1992));
   NAND2_X1 i_2256 (.A1(A[23]), .A2(B[11]), .ZN(n_2003));
   NOR2_X1 i_2257 (.A1(n_2003), .A2(n_1954), .ZN(n_2025));
   AOI22_X1 i_2258 (.A1(A[23]), .A2(B[9]), .B1(A[21]), .B2(B[11]), .ZN(n_2026));
   NOR2_X1 i_2259 (.A1(n_2025), .A2(n_2026), .ZN(n_2037));
   XNOR2_X1 i_2260 (.A(n_2037), .B(n_1992), .ZN(n_2038));
   INV_X1 i_2261 (.A(n_1933), .ZN(n_2039));
   INV_X1 i_2262 (.A(n_1932), .ZN(n_2040));
   OAI22_X1 i_2263 (.A1(n_2039), .A2(n_1934), .B1(n_2040), .B2(n_1726), .ZN(
      n_2041));
   INV_X1 i_2264 (.A(n_2041), .ZN(n_2052));
   AOI22_X1 i_2265 (.A1(n_1850), .A2(n_1853), .B1(n_1849), .B2(n_1843), .ZN(
      n_2053));
   NOR2_X1 i_2266 (.A1(n_1992), .A2(n_1954), .ZN(n_2054));
   AOI22_X1 i_2267 (.A1(B[10]), .A2(A[21]), .B1(B[9]), .B2(A[22]), .ZN(n_2055));
   NOR2_X1 i_2268 (.A1(n_2054), .A2(n_2055), .ZN(n_2056));
   AND2_X1 i_2269 (.A1(B[11]), .A2(A[20]), .ZN(n_2057));
   XOR2_X1 i_2270 (.A(n_2056), .B(n_2057), .Z(n_2058));
   XNOR2_X1 i_2271 (.A(n_2053), .B(n_2041), .ZN(n_2059));
   NAND2_X1 i_2272 (.A1(n_2058), .A2(n_2059), .ZN(n_2060));
   OAI21_X1 i_2273 (.A(n_2060), .B1(n_2059), .B2(n_2058), .ZN(n_2061));
   AOI22_X1 i_2274 (.A1(n_1842), .A2(n_1833), .B1(n_1832), .B2(n_1813), .ZN(
      n_2062));
   NAND2_X1 i_2275 (.A1(n_2061), .A2(n_2062), .ZN(n_2063));
   OAI21_X1 i_2276 (.A(n_2063), .B1(n_2062), .B2(n_2061), .ZN(n_2064));
   INV_X1 i_2277 (.A(n_1795), .ZN(n_2065));
   AOI22_X1 i_2278 (.A1(n_2065), .A2(n_1796), .B1(n_1811), .B2(n_1797), .ZN(
      n_2066));
   INV_X1 i_2279 (.A(n_2066), .ZN(n_2067));
   OAI21_X1 i_2280 (.A(n_2063), .B1(n_2064), .B2(n_2067), .ZN(n_2068));
   XNOR2_X1 i_2281 (.A(n_1976), .B(n_1981), .ZN(n_2069));
   XOR2_X1 i_2282 (.A(n_1991), .B(n_2038), .Z(n_2070));
   XOR2_X1 i_2283 (.A(n_2069), .B(n_2070), .Z(n_2071));
   INV_X1 i_2284 (.A(n_2068), .ZN(n_2072));
   AOI22_X1 i_2285 (.A1(n_2071), .A2(n_2072), .B1(n_2069), .B2(n_2070), .ZN(
      n_2073));
   XNOR2_X1 i_2286 (.A(n_2133), .B(n_2075), .ZN(n_2074));
   AOI21_X1 i_2287 (.A(n_2077), .B1(n_2085), .B2(n_2076), .ZN(n_2075));
   AOI21_X1 i_2288 (.A(n_2077), .B1(n_2079), .B2(n_2078), .ZN(n_2076));
   NOR2_X1 i_2289 (.A1(n_2079), .A2(n_2078), .ZN(n_2077));
   AOI21_X1 i_2290 (.A(n_2082), .B1(n_2081), .B2(n_2080), .ZN(n_2078));
   XOR2_X1 i_2291 (.A(n_2003), .B(n_2149), .Z(n_2079));
   XNOR2_X1 i_2292 (.A(n_2175), .B(n_2174), .ZN(n_2080));
   AOI21_X1 i_2293 (.A(n_2082), .B1(n_2084), .B2(n_2083), .ZN(n_2081));
   NOR2_X1 i_2294 (.A1(n_2084), .A2(n_2083), .ZN(n_2082));
   XOR2_X1 i_2295 (.A(n_2153), .B(n_2152), .Z(n_2083));
   XOR2_X1 i_2296 (.A(n_1958), .B(n_2200), .Z(n_2084));
   AOI21_X1 i_2297 (.A(n_2114), .B1(n_2111), .B2(n_2086), .ZN(n_2085));
   OAI22_X1 i_2298 (.A1(n_2107), .A2(n_2088), .B1(n_2108), .B2(n_2087), .ZN(
      n_2086));
   INV_X1 i_2299 (.A(n_2088), .ZN(n_2087));
   NAND2_X1 i_2300 (.A1(B[11]), .A2(A[22]), .ZN(n_2088));
   INV_X1 i_2301 (.A(n_2108), .ZN(n_2107));
   XOR2_X1 i_2302 (.A(n_2110), .B(n_2109), .Z(n_2108));
   NOR2_X1 i_2303 (.A1(n_2243), .A2(n_1792), .ZN(n_2109));
   AOI21_X1 i_2304 (.A(n_2025), .B1(n_2236), .B2(n_2037), .ZN(n_2110));
   AOI21_X1 i_2305 (.A(n_2114), .B1(n_2116), .B2(n_2115), .ZN(n_2111));
   NOR2_X1 i_2306 (.A1(n_2116), .A2(n_2115), .ZN(n_2114));
   AOI21_X1 i_2307 (.A(n_2126), .B1(n_2125), .B2(n_2118), .ZN(n_2115));
   INV_X1 i_2308 (.A(n_2117), .ZN(n_2116));
   OAI33_X1 i_2309 (.A1(n_1235), .A2(n_1368), .A3(n_2132), .B1(n_1979), .B2(
      n_339), .B3(n_1533), .ZN(n_2117));
   OAI21_X1 i_2310 (.A(n_2124), .B1(n_1964), .B2(n_2119), .ZN(n_2118));
   NAND2_X1 i_2311 (.A1(n_2124), .A2(n_2122), .ZN(n_2119));
   INV_X1 i_2312 (.A(n_2123), .ZN(n_2122));
   AOI22_X1 i_2313 (.A1(B[16]), .A2(A[15]), .B1(B[17]), .B2(A[14]), .ZN(n_2123));
   OR2_X1 i_2314 (.A1(n_1963), .A2(n_1848), .ZN(n_2124));
   AOI21_X1 i_2315 (.A(n_2126), .B1(n_2129), .B2(n_2127), .ZN(n_2125));
   NOR2_X1 i_2316 (.A1(n_2129), .A2(n_2127), .ZN(n_2126));
   INV_X1 i_2317 (.A(n_2128), .ZN(n_2127));
   OAI22_X1 i_2318 (.A1(n_1924), .A2(n_2234), .B1(n_2131), .B2(n_2130), .ZN(
      n_2128));
   AOI21_X1 i_2319 (.A(n_2054), .B1(n_2056), .B2(n_2057), .ZN(n_2129));
   NAND2_X1 i_2320 (.A1(B[14]), .A2(A[17]), .ZN(n_2130));
   XNOR2_X1 i_2321 (.A(n_1924), .B(n_2234), .ZN(n_2131));
   NAND2_X1 i_2322 (.A1(B[21]), .A2(A[10]), .ZN(n_2132));
   XNOR2_X1 i_2323 (.A(n_2178), .B(n_2134), .ZN(n_2133));
   XOR2_X1 i_2324 (.A(n_2146), .B(n_2135), .Z(n_2134));
   XOR2_X1 i_2325 (.A(n_2137), .B(n_2136), .Z(n_2135));
   NOR2_X1 i_2326 (.A1(n_229), .A2(n_1881), .ZN(n_2136));
   NOR2_X1 i_2327 (.A1(n_2143), .A2(n_2142), .ZN(n_2137));
   AOI22_X1 i_2328 (.A1(B[12]), .A2(A[23]), .B1(B[14]), .B2(A[21]), .ZN(n_2142));
   AND3_X1 i_2329 (.A1(B[12]), .A2(A[21]), .A3(n_2145), .ZN(n_2143));
   NOR2_X1 i_2330 (.A1(n_559), .A2(n_1792), .ZN(n_2145));
   XOR2_X1 i_2331 (.A(n_2148), .B(n_2147), .Z(n_2146));
   OAI22_X1 i_2332 (.A1(n_2215), .A2(n_2184), .B1(n_2183), .B2(n_2182), .ZN(
      n_2147));
   OAI21_X1 i_2333 (.A(n_2150), .B1(n_2003), .B2(n_2149), .ZN(n_2148));
   OAI21_X1 i_2334 (.A(n_2150), .B1(n_2173), .B2(n_2151), .ZN(n_2149));
   NAND2_X1 i_2335 (.A1(n_2173), .A2(n_2151), .ZN(n_2150));
   OAI22_X1 i_2336 (.A1(n_1985), .A2(n_2177), .B1(n_2153), .B2(n_2152), .ZN(
      n_2151));
   OR2_X1 i_2337 (.A1(n_559), .A2(n_853), .ZN(n_2152));
   OAI21_X1 i_2338 (.A(n_2154), .B1(n_1985), .B2(n_2177), .ZN(n_2153));
   INV_X1 i_2339 (.A(n_2172), .ZN(n_2154));
   AOI22_X1 i_2340 (.A1(B[13]), .A2(A[20]), .B1(B[12]), .B2(A[21]), .ZN(n_2172));
   OAI22_X1 i_2341 (.A1(n_1965), .A2(n_2176), .B1(n_2175), .B2(n_2174), .ZN(
      n_2173));
   NAND2_X1 i_2342 (.A1(B[15]), .A2(A[18]), .ZN(n_2174));
   XNOR2_X1 i_2343 (.A(n_1965), .B(n_2176), .ZN(n_2175));
   NAND2_X1 i_2344 (.A1(B[17]), .A2(A[16]), .ZN(n_2176));
   NAND2_X1 i_2345 (.A1(B[13]), .A2(A[21]), .ZN(n_2177));
   AOI22_X1 i_2346 (.A1(n_2181), .A2(n_2180), .B1(n_2194), .B2(n_2179), .ZN(
      n_2178));
   XOR2_X1 i_2347 (.A(n_2181), .B(n_2180), .Z(n_2179));
   XOR2_X1 i_2348 (.A(n_2186), .B(n_2185), .Z(n_2180));
   XOR2_X1 i_2349 (.A(n_2183), .B(n_2182), .Z(n_2181));
   NAND2_X1 i_2350 (.A1(B[23]), .A2(A[11]), .ZN(n_2182));
   XNOR2_X1 i_2351 (.A(n_2215), .B(n_2184), .ZN(n_2183));
   NAND2_X1 i_2352 (.A1(B[21]), .A2(A[13]), .ZN(n_2184));
   NOR2_X1 i_2353 (.A1(n_557), .A2(n_856), .ZN(n_2185));
   AOI21_X1 i_2354 (.A(n_2188), .B1(n_2209), .B2(n_2187), .ZN(n_2186));
   NAND2_X1 i_2355 (.A1(B[18]), .A2(A[16]), .ZN(n_2187));
   NOR3_X1 i_2356 (.A1(n_1305), .A2(n_2209), .A3(n_1532), .ZN(n_2188));
   XNOR2_X1 i_2357 (.A(n_2216), .B(n_2195), .ZN(n_2194));
   XOR2_X1 i_2358 (.A(n_2210), .B(n_2199), .Z(n_2195));
   INV_X1 i_2359 (.A(n_2199), .ZN(n_2196));
   OAI22_X1 i_2360 (.A1(n_1957), .A2(n_2209), .B1(n_1958), .B2(n_2200), .ZN(
      n_2199));
   OAI21_X1 i_2361 (.A(n_2201), .B1(n_1957), .B2(n_2209), .ZN(n_2200));
   INV_X1 i_2362 (.A(n_2202), .ZN(n_2201));
   AOI22_X1 i_2363 (.A1(B[19]), .A2(A[14]), .B1(B[18]), .B2(A[15]), .ZN(n_2202));
   NAND2_X1 i_2364 (.A1(B[19]), .A2(A[15]), .ZN(n_2209));
   OAI22_X1 i_2365 (.A1(n_1977), .A2(n_2215), .B1(n_2212), .B2(n_2211), .ZN(
      n_2210));
   NAND2_X1 i_2366 (.A1(B[23]), .A2(A[10]), .ZN(n_2211));
   OAI21_X1 i_2367 (.A(n_2213), .B1(n_1977), .B2(n_2215), .ZN(n_2212));
   INV_X1 i_2368 (.A(n_2214), .ZN(n_2213));
   AOI22_X1 i_2369 (.A1(B[22]), .A2(A[11]), .B1(B[21]), .B2(A[12]), .ZN(n_2214));
   NAND2_X1 i_2370 (.A1(B[22]), .A2(A[12]), .ZN(n_2215));
   AOI22_X1 i_2371 (.A1(n_2235), .A2(n_2233), .B1(n_2218), .B2(n_2217), .ZN(
      n_2216));
   AOI21_X1 i_2372 (.A(n_1960), .B1(n_2242), .B2(n_1957), .ZN(n_2217));
   XOR2_X1 i_2373 (.A(n_2235), .B(n_2233), .Z(n_2218));
   OAI33_X1 i_2374 (.A1(n_229), .A2(n_1322), .A3(n_2234), .B1(n_1987), .B2(n_559), 
      .B3(n_1028), .ZN(n_2233));
   NAND2_X1 i_2375 (.A1(B[12]), .A2(A[19]), .ZN(n_2234));
   OAI21_X1 i_2376 (.A(n_2244), .B1(n_1967), .B2(n_1963), .ZN(n_2235));
   INV_X1 i_2377 (.A(n_1992), .ZN(n_2236));
   INV_X1 i_2378 (.A(n_1959), .ZN(n_2242));
   INV_X1 i_2379 (.A(B[10]), .ZN(n_2243));
   INV_X1 i_2380 (.A(n_1966), .ZN(n_2244));
   NAND2_X1 i_2381 (.A1(B[12]), .A2(A[22]), .ZN(n_2245));
   XNOR2_X1 i_2382 (.A(n_2245), .B(n_2177), .ZN(n_2246));
   NAND2_X1 i_2383 (.A1(A[20]), .A2(B[14]), .ZN(n_2248));
   NAND2_X1 i_2384 (.A1(B[15]), .A2(A[19]), .ZN(n_2249));
   AND2_X1 i_2385 (.A1(A[18]), .A2(B[16]), .ZN(n_2250));
   INV_X1 i_2387 (.A(n_2249), .ZN(n_2251));
   NAND2_X1 i_2388 (.A1(n_2250), .A2(n_2251), .ZN(n_2252));
   OAI21_X1 i_2389 (.A(n_2252), .B1(n_2251), .B2(n_2250), .ZN(n_2253));
   NAND2_X1 i_2390 (.A1(A[17]), .A2(B[17]), .ZN(n_2256));
   OAI21_X1 i_2391 (.A(n_2252), .B1(n_2253), .B2(n_2256), .ZN(n_2257));
   OAI22_X1 i_2392 (.A1(n_2246), .A2(n_2248), .B1(n_2245), .B2(n_2177), .ZN(
      n_2258));
   NAND2_X1 i_2393 (.A1(n_2257), .A2(n_2258), .ZN(n_2259));
   OAI21_X1 i_2394 (.A(n_2259), .B1(n_2258), .B2(n_2257), .ZN(n_2260));
   AOI21_X1 i_2395 (.A(n_2188), .B1(n_2186), .B2(n_2185), .ZN(n_2261));
   NAND2_X1 i_2396 (.A1(B[16]), .A2(A[20]), .ZN(n_2266));
   NAND2_X1 i_2397 (.A1(B[15]), .A2(A[21]), .ZN(n_2267));
   NOR2_X1 i_2398 (.A1(n_2266), .A2(n_2267), .ZN(n_2268));
   INV_X1 i_2399 (.A(n_2268), .ZN(n_2269));
   AOI21_X1 i_2400 (.A(n_2268), .B1(n_2266), .B2(n_2267), .ZN(n_2270));
   INV_X1 i_2401 (.A(n_2270), .ZN(n_2271));
   NAND2_X1 i_2402 (.A1(B[17]), .A2(A[19]), .ZN(n_2272));
   OAI21_X1 i_2403 (.A(n_2259), .B1(n_2260), .B2(n_2261), .ZN(n_2273));
   XNOR2_X1 i_2404 (.A(n_2270), .B(n_2272), .ZN(n_2274));
   NOR2_X1 i_2405 (.A1(n_2273), .A2(n_2274), .ZN(n_2275));
   AOI21_X1 i_2406 (.A(n_2143), .B1(n_2137), .B2(n_2136), .ZN(n_2276));
   NAND2_X1 i_2407 (.A1(B[13]), .A2(A[23]), .ZN(n_2277));
   NAND2_X1 i_2408 (.A1(B[14]), .A2(A[22]), .ZN(n_2278));
   XNOR2_X1 i_2409 (.A(n_2276), .B(n_2277), .ZN(n_2279));
   XNOR2_X1 i_2410 (.A(n_2279), .B(n_2278), .ZN(n_2280));
   NAND2_X1 i_2411 (.A1(n_2273), .A2(n_2274), .ZN(n_2281));
   AOI21_X1 i_2412 (.A(n_2275), .B1(n_2281), .B2(n_2280), .ZN(n_2302));
   INV_X1 i_2413 (.A(n_2302), .ZN(n_2303));
   INV_X1 i_2414 (.A(n_2305), .ZN(n_2304));
   AOI21_X1 i_2415 (.A(n_2307), .B1(n_2322), .B2(n_2306), .ZN(n_2305));
   AOI21_X1 i_2416 (.A(n_2307), .B1(n_2310), .B2(n_2308), .ZN(n_2306));
   NOR2_X1 i_2417 (.A1(n_2310), .A2(n_2308), .ZN(n_2307));
   INV_X1 i_2418 (.A(n_2309), .ZN(n_2308));
   OAI22_X1 i_2419 (.A1(n_2355), .A2(n_2320), .B1(n_2319), .B2(n_2318), .ZN(
      n_2309));
   AOI21_X1 i_2420 (.A(n_2316), .B1(n_2312), .B2(n_2311), .ZN(n_2310));
   NOR2_X1 i_2421 (.A1(n_558), .A2(n_1533), .ZN(n_2311));
   NOR2_X1 i_2422 (.A1(n_2316), .A2(n_2314), .ZN(n_2312));
   AOI22_X1 i_2423 (.A1(A[16]), .A2(B[22]), .B1(A[17]), .B2(B[21]), .ZN(n_2314));
   NOR2_X1 i_2424 (.A1(n_2327), .A2(n_2317), .ZN(n_2316));
   NAND2_X1 i_2425 (.A1(A[17]), .A2(B[22]), .ZN(n_2317));
   NAND2_X1 i_2426 (.A1(A[18]), .A2(B[20]), .ZN(n_2318));
   XNOR2_X1 i_2427 (.A(n_2355), .B(n_2320), .ZN(n_2319));
   NAND2_X1 i_2428 (.A1(A[20]), .A2(B[18]), .ZN(n_2320));
   OAI21_X1 i_2429 (.A(n_2331), .B1(n_2330), .B2(n_2323), .ZN(n_2322));
   INV_X1 i_2430 (.A(n_2324), .ZN(n_2323));
   OAI22_X1 i_2432 (.A1(n_2329), .A2(n_2327), .B1(n_2326), .B2(n_2325), .ZN(
      n_2324));
   NAND2_X1 i_2433 (.A1(A[14]), .A2(B[23]), .ZN(n_2325));
   XNOR2_X1 i_2434 (.A(n_2329), .B(n_2327), .ZN(n_2326));
   NAND2_X1 i_2435 (.A1(A[16]), .A2(B[21]), .ZN(n_2327));
   NAND2_X1 i_2436 (.A1(A[15]), .A2(B[22]), .ZN(n_2329));
   OAI21_X1 i_2437 (.A(n_2331), .B1(n_2333), .B2(n_2332), .ZN(n_2330));
   NAND2_X1 i_2438 (.A1(n_2333), .A2(n_2332), .ZN(n_2331));
   OAI22_X1 i_2439 (.A1(n_2267), .A2(n_2339), .B1(n_2336), .B2(n_2335), .ZN(
      n_2332));
   OAI22_X1 i_2440 (.A1(n_2356), .A2(n_2355), .B1(n_2341), .B2(n_2340), .ZN(
      n_2333));
   NAND2_X1 i_2441 (.A1(A[20]), .A2(B[17]), .ZN(n_2335));
   OAI21_X1 i_2442 (.A(n_2337), .B1(n_2267), .B2(n_2339), .ZN(n_2336));
   INV_X1 i_2443 (.A(n_2338), .ZN(n_2337));
   AOI22_X1 i_2444 (.A1(A[22]), .A2(B[15]), .B1(A[21]), .B2(B[16]), .ZN(n_2338));
   NAND2_X1 i_2445 (.A1(A[22]), .A2(B[16]), .ZN(n_2339));
   NAND2_X1 i_2446 (.A1(A[17]), .A2(B[20]), .ZN(n_2340));
   OAI21_X1 i_2447 (.A(n_2353), .B1(n_2356), .B2(n_2355), .ZN(n_2341));
   INV_X1 i_2448 (.A(n_2354), .ZN(n_2353));
   AOI22_X1 i_2449 (.A1(A[18]), .A2(B[19]), .B1(A[19]), .B2(B[18]), .ZN(n_2354));
   NAND2_X1 i_2450 (.A1(A[19]), .A2(B[19]), .ZN(n_2355));
   NAND2_X1 i_2451 (.A1(A[18]), .A2(B[18]), .ZN(n_2356));
   XOR2_X1 i_2452 (.A(n_2371), .B(n_2360), .Z(n_2357));
   OAI22_X1 i_2453 (.A1(n_2317), .A2(n_2370), .B1(n_2363), .B2(n_2361), .ZN(
      n_2360));
   NAND2_X1 i_2454 (.A1(B[21]), .A2(A[19]), .ZN(n_2361));
   NOR2_X1 i_2455 (.A1(n_2364), .A2(n_2363), .ZN(n_2362));
   AOI22_X1 i_2456 (.A1(B[23]), .A2(A[17]), .B1(B[22]), .B2(A[18]), .ZN(n_2363));
   NOR2_X1 i_2457 (.A1(n_2317), .A2(n_2370), .ZN(n_2364));
   NAND2_X1 i_2458 (.A1(B[23]), .A2(A[18]), .ZN(n_2370));
   INV_X1 i_2459 (.A(n_2372), .ZN(n_2371));
   AOI21_X1 i_2460 (.A(n_2377), .B1(n_2374), .B2(n_2373), .ZN(n_2372));
   NOR2_X1 i_2461 (.A1(n_1322), .A2(n_856), .ZN(n_2373));
   NOR2_X1 i_2462 (.A1(n_2377), .A2(n_2376), .ZN(n_2374));
   AOI22_X1 i_2463 (.A1(B[19]), .A2(A[21]), .B1(B[18]), .B2(A[22]), .ZN(n_2376));
   NOR2_X1 i_2464 (.A1(n_2381), .A2(n_2378), .ZN(n_2377));
   NAND2_X1 i_2465 (.A1(B[19]), .A2(A[22]), .ZN(n_2378));
   NAND2_X1 i_2466 (.A1(B[18]), .A2(A[21]), .ZN(n_2381));
   XOR2_X1 i_2467 (.A(n_2405), .B(n_2383), .Z(n_2382));
   XOR2_X1 i_2468 (.A(n_2400), .B(n_2384), .Z(n_2383));
   XNOR2_X1 i_2469 (.A(n_2362), .B(n_2361), .ZN(n_2384));
   XOR2_X1 i_2470 (.A(n_2404), .B(n_2403), .Z(n_2400));
   OAI22_X1 i_2471 (.A1(n_2339), .A2(n_2430), .B1(n_2410), .B2(n_2408), .ZN(
      n_2403));
   XOR2_X1 i_2472 (.A(n_2374), .B(n_2373), .Z(n_2404));
   XNOR2_X1 i_2473 (.A(n_2420), .B(n_2406), .ZN(n_2405));
   AOI22_X1 i_2474 (.A1(n_2419), .A2(n_2418), .B1(n_2417), .B2(n_2407), .ZN(
      n_2406));
   XOR2_X1 i_2475 (.A(n_2410), .B(n_2408), .Z(n_2407));
   OAI21_X1 i_2476 (.A(n_2409), .B1(n_2339), .B2(n_2430), .ZN(n_2408));
   OAI22_X1 i_2480 (.A1(n_1232), .A2(n_1881), .B1(n_592), .B2(n_1792), .ZN(
      n_2409));
   AOI21_X1 i_2481 (.A(n_2413), .B1(n_2443), .B2(n_2411), .ZN(n_2410));
   NOR2_X1 i_2482 (.A1(n_2413), .A2(n_2412), .ZN(n_2411));
   AOI22_X1 i_2483 (.A1(A[23]), .A2(B[15]), .B1(A[21]), .B2(B[17]), .ZN(n_2412));
   NOR2_X1 i_2484 (.A1(n_2267), .A2(n_2430), .ZN(n_2413));
   XOR2_X1 i_2485 (.A(n_2419), .B(n_2418), .Z(n_2417));
   XOR2_X1 i_2486 (.A(n_2425), .B(n_2424), .Z(n_2418));
   XOR2_X1 i_2487 (.A(n_2433), .B(n_2432), .Z(n_2419));
   XNOR2_X1 i_2488 (.A(n_2305), .B(n_2421), .ZN(n_2420));
   XOR2_X1 i_2489 (.A(n_2423), .B(n_2422), .Z(n_2421));
   AOI21_X1 i_2490 (.A(n_2428), .B1(n_2431), .B2(n_2429), .ZN(n_2422));
   OAI22_X1 i_2491 (.A1(n_2381), .A2(n_2426), .B1(n_2425), .B2(n_2424), .ZN(
      n_2423));
   NAND2_X1 i_2492 (.A1(A[19]), .A2(B[20]), .ZN(n_2424));
   XNOR2_X1 i_2493 (.A(n_2381), .B(n_2426), .ZN(n_2425));
   NAND2_X1 i_2494 (.A1(A[20]), .A2(B[19]), .ZN(n_2426));
   NAND2_X1 i_2495 (.A1(n_2431), .A2(n_2429), .ZN(n_2427));
   NOR2_X1 i_2496 (.A1(n_2431), .A2(n_2429), .ZN(n_2428));
   INV_X1 i_2497 (.A(n_2430), .ZN(n_2429));
   NAND2_X1 i_2498 (.A1(A[23]), .A2(B[17]), .ZN(n_2430));
   OAI22_X1 i_2499 (.A1(n_2317), .A2(n_2442), .B1(n_2433), .B2(n_2432), .ZN(
      n_2431));
   NAND2_X1 i_2500 (.A1(A[16]), .A2(B[23]), .ZN(n_2432));
   XNOR2_X1 i_2501 (.A(n_2317), .B(n_2442), .ZN(n_2433));
   NAND2_X1 i_2502 (.A1(A[18]), .A2(B[21]), .ZN(n_2442));
   INV_X1 i_2503 (.A(n_2339), .ZN(n_2443));
   AOI21_X1 i_2504 (.A(n_2446), .B1(n_2460), .B2(n_2445), .ZN(n_2444));
   AOI21_X1 i_2505 (.A(n_2446), .B1(n_2448), .B2(n_2447), .ZN(n_2445));
   NOR2_X1 i_2506 (.A1(n_2448), .A2(n_2447), .ZN(n_2446));
   XOR2_X1 i_2507 (.A(n_2322), .B(n_2306), .Z(n_2447));
   AOI22_X1 i_2508 (.A1(n_2453), .A2(n_2451), .B1(n_2450), .B2(n_2449), .ZN(
      n_2448));
   XOR2_X1 i_2509 (.A(n_2411), .B(n_2339), .Z(n_2449));
   XOR2_X1 i_2510 (.A(n_2453), .B(n_2451), .Z(n_2450));
   XNOR2_X1 i_2511 (.A(n_2319), .B(n_2318), .ZN(n_2451));
   AOI22_X1 i_2512 (.A1(n_2145), .A2(n_2456), .B1(n_2455), .B2(n_2454), .ZN(
      n_2453));
   OAI21_X1 i_2513 (.A(n_2269), .B1(n_2271), .B2(n_2272), .ZN(n_2454));
   XOR2_X1 i_2514 (.A(n_2145), .B(n_2456), .Z(n_2455));
   OAI21_X1 i_2516 (.A(n_2457), .B1(n_2340), .B2(n_2505), .ZN(n_2456));
   NAND2_X1 i_2517 (.A1(n_2506), .A2(n_2458), .ZN(n_2457));
   AOI21_X1 i_2518 (.A(n_2459), .B1(n_2507), .B2(n_2504), .ZN(n_2458));
   AOI22_X1 i_2519 (.A1(A[17]), .A2(B[19]), .B1(A[16]), .B2(B[20]), .ZN(n_2459));
   AOI21_X1 i_2520 (.A(n_2463), .B1(n_2462), .B2(n_2461), .ZN(n_2460));
   XNOR2_X1 i_2521 (.A(n_2330), .B(n_2324), .ZN(n_2461));
   AOI21_X1 i_2522 (.A(n_2463), .B1(n_2465), .B2(n_2464), .ZN(n_2462));
   NOR2_X1 i_2523 (.A1(n_2465), .A2(n_2464), .ZN(n_2463));
   XNOR2_X1 i_2524 (.A(n_2312), .B(n_2311), .ZN(n_2464));
   AOI21_X1 i_2525 (.A(n_2468), .B1(n_2467), .B2(n_2466), .ZN(n_2465));
   OAI22_X1 i_2526 (.A1(n_2279), .A2(n_2278), .B1(n_2276), .B2(n_2277), .ZN(
      n_2466));
   AOI21_X1 i_2527 (.A(n_2468), .B1(n_2479), .B2(n_2469), .ZN(n_2467));
   NOR2_X1 i_2528 (.A1(n_2479), .A2(n_2469), .ZN(n_2468));
   OAI22_X1 i_2529 (.A1(n_2494), .A2(n_2493), .B1(n_2491), .B2(n_2484), .ZN(
      n_2469));
   AOI21_X1 i_2530 (.A(n_2483), .B1(n_2481), .B2(n_2480), .ZN(n_2479));
   NOR2_X1 i_2531 (.A1(n_256), .A2(n_1533), .ZN(n_2480));
   NOR2_X1 i_2532 (.A1(n_2483), .A2(n_2482), .ZN(n_2481));
   AOI22_X1 i_2533 (.A1(A[14]), .A2(B[22]), .B1(A[15]), .B2(B[21]), .ZN(n_2482));
   NOR3_X1 i_2534 (.A1(n_2516), .A2(n_2508), .A3(n_2329), .ZN(n_2483));
   OAI21_X1 i_2535 (.A(n_2487), .B1(n_2486), .B2(n_2485), .ZN(n_2484));
   NAND2_X1 i_2536 (.A1(A[12]), .A2(B[23]), .ZN(n_2485));
   OAI21_X1 i_2537 (.A(n_2487), .B1(n_2489), .B2(n_2488), .ZN(n_2486));
   NAND2_X1 i_2538 (.A1(n_2489), .A2(n_2488), .ZN(n_2487));
   NOR2_X1 i_2539 (.A1(n_256), .A2(n_1368), .ZN(n_2488));
   NOR2_X1 i_2540 (.A1(n_2516), .A2(n_2508), .ZN(n_2489));
   OAI21_X1 i_2541 (.A(n_2492), .B1(n_2494), .B2(n_2493), .ZN(n_2490));
   INV_X1 i_2542 (.A(n_2492), .ZN(n_2491));
   NAND2_X1 i_2543 (.A1(n_2494), .A2(n_2493), .ZN(n_2492));
   OAI21_X1 i_2544 (.A(n_2502), .B1(n_2501), .B2(n_2500), .ZN(n_2493));
   OAI21_X1 i_2545 (.A(n_2499), .B1(n_2496), .B2(n_2495), .ZN(n_2494));
   NAND2_X1 i_2546 (.A1(A[18]), .A2(B[17]), .ZN(n_2495));
   NAND2_X1 i_2547 (.A1(n_2499), .A2(n_2497), .ZN(n_2496));
   INV_X1 i_2548 (.A(n_2498), .ZN(n_2497));
   AOI22_X1 i_2549 (.A1(A[19]), .A2(B[16]), .B1(A[20]), .B2(B[15]), .ZN(n_2498));
   OR2_X1 i_2550 (.A1(n_2249), .A2(n_2266), .ZN(n_2499));
   NAND2_X1 i_2552 (.A1(A[17]), .A2(B[18]), .ZN(n_2500));
   OAI21_X1 i_2553 (.A(n_2502), .B1(n_2504), .B2(n_2503), .ZN(n_2501));
   NAND2_X1 i_2554 (.A1(n_2504), .A2(n_2503), .ZN(n_2502));
   NOR2_X1 i_2555 (.A1(n_558), .A2(n_856), .ZN(n_2503));
   INV_X1 i_2556 (.A(n_2505), .ZN(n_2504));
   NAND2_X1 i_2557 (.A1(A[16]), .A2(B[19]), .ZN(n_2505));
   INV_X1 i_2558 (.A(n_2356), .ZN(n_2506));
   INV_X1 i_2559 (.A(n_2340), .ZN(n_2507));
   INV_X1 i_2560 (.A(B[21]), .ZN(n_2508));
   INV_X1 i_2561 (.A(A[14]), .ZN(n_2516));
   NAND2_X1 i_2562 (.A1(A[22]), .A2(B[22]), .ZN(n_2517));
   NOR2_X1 i_2563 (.A1(n_1322), .A2(n_1533), .ZN(n_2518));
   NAND2_X1 i_2564 (.A1(A[21]), .A2(B[23]), .ZN(n_2519));
   XNOR2_X1 i_2565 (.A(n_2517), .B(n_2519), .ZN(n_2520));
   INV_X1 i_2566 (.A(n_2378), .ZN(n_2521));
   NAND2_X1 i_2567 (.A1(B[20]), .A2(A[23]), .ZN(n_2523));
   NOR2_X1 i_2568 (.A1(n_2523), .A2(n_2381), .ZN(n_2524));
   AOI22_X1 i_2569 (.A1(A[21]), .A2(B[20]), .B1(B[18]), .B2(A[23]), .ZN(n_2525));
   NOR2_X1 i_2570 (.A1(n_2524), .A2(n_2525), .ZN(n_2526));
   NAND2_X1 i_2571 (.A1(n_2526), .A2(n_2521), .ZN(n_2528));
   INV_X1 i_2572 (.A(n_2524), .ZN(n_2529));
   NAND2_X1 i_2573 (.A1(n_2528), .A2(n_2529), .ZN(n_2530));
   AOI21_X1 i_2574 (.A(n_2530), .B1(B[19]), .B2(A[23]), .ZN(n_2531));
   NAND2_X1 i_2575 (.A1(B[20]), .A2(A[22]), .ZN(n_2532));
   NAND3_X1 i_2576 (.A1(n_2530), .A2(B[19]), .A3(A[23]), .ZN(n_2533));
   NAND2_X1 i_2577 (.A1(B[22]), .A2(A[20]), .ZN(n_2541));
   NAND2_X1 i_2578 (.A1(B[21]), .A2(A[21]), .ZN(n_2554));
   XNOR2_X1 i_2579 (.A(n_2554), .B(n_2541), .ZN(n_2555));
   NAND2_X1 i_2580 (.A1(B[23]), .A2(A[19]), .ZN(n_2556));
   AOI21_X1 i_2581 (.A(n_2531), .B1(n_2532), .B2(n_2533), .ZN(n_2557));
   OAI22_X1 i_2582 (.A1(n_2555), .A2(n_2556), .B1(n_2554), .B2(n_2541), .ZN(
      n_2558));
   XOR2_X1 i_2583 (.A(n_2557), .B(n_2558), .Z(n_2559));
   INV_X1 i_2584 (.A(n_2523), .ZN(n_2560));
   AOI22_X1 i_2585 (.A1(n_2559), .A2(n_2560), .B1(n_2557), .B2(n_2558), .ZN(
      n_2561));
   NAND2_X1 i_2586 (.A1(B[21]), .A2(A[23]), .ZN(n_2562));
   XNOR2_X1 i_2590 (.A(n_2520), .B(n_2562), .ZN(n_2563));
   AOI22_X1 i_2596 (.A1(A[21]), .A2(B[22]), .B1(B[21]), .B2(A[22]), .ZN(n_2564));
   INV_X1 i_2597 (.A(n_2564), .ZN(n_2565));
   NOR2_X1 i_2598 (.A1(n_2554), .A2(n_2517), .ZN(n_2566));
   OAI21_X1 i_2599 (.A(n_2565), .B1(n_2566), .B2(n_2518), .ZN(n_2567));
   XOR2_X1 i_2600 (.A(n_2563), .B(n_2567), .Z(n_2568));
   AOI22_X1 i_2601 (.A1(n_2561), .A2(n_2568), .B1(n_2563), .B2(n_2567), .ZN(
      n_2569));
   INV_X1 i_2602 (.A(n_2569), .ZN(n_2570));
   NOR2_X1 i_2603 (.A1(n_2566), .A2(n_2564), .ZN(n_2571));
   NAND2_X1 i_2604 (.A1(n_2582), .A2(n_2581), .ZN(n_2580));
   XNOR2_X1 i_2605 (.A(n_2561), .B(n_2568), .ZN(n_2581));
   OAI21_X1 i_2606 (.A(n_2593), .B1(n_2592), .B2(n_2583), .ZN(n_2582));
   AOI22_X1 i_2607 (.A1(n_2586), .A2(n_2585), .B1(n_2590), .B2(n_2584), .ZN(
      n_2583));
   XOR2_X1 i_2608 (.A(n_2586), .B(n_2585), .Z(n_2584));
   XOR2_X1 i_2609 (.A(n_2555), .B(n_2556), .Z(n_2585));
   OAI22_X1 i_2610 (.A1(n_2361), .A2(n_2541), .B1(n_2370), .B2(n_2588), .ZN(
      n_2586));
   NOR2_X1 i_2611 (.A1(n_2589), .A2(n_2588), .ZN(n_2587));
   AOI22_X1 i_2612 (.A1(A[20]), .A2(B[21]), .B1(A[19]), .B2(B[22]), .ZN(n_2588));
   NOR2_X1 i_2613 (.A1(n_2361), .A2(n_2541), .ZN(n_2589));
   XNOR2_X1 i_2623 (.A(n_2532), .B(n_2591), .ZN(n_2590));
   NOR2_X1 i_2624 (.A1(n_2531), .A2(n_2600), .ZN(n_2591));
   OAI21_X1 i_2625 (.A(n_2593), .B1(n_2599), .B2(n_2598), .ZN(n_2592));
   NAND2_X1 i_2626 (.A1(n_2599), .A2(n_2598), .ZN(n_2593));
   XOR2_X1 i_2627 (.A(n_2571), .B(n_2518), .Z(n_2598));
   XNOR2_X1 i_2628 (.A(n_2559), .B(n_2523), .ZN(n_2599));
   INV_X1 i_2629 (.A(n_2533), .ZN(n_2600));
endmodule

module N_Bit_Mult(A, B, Out);
   input [23:0]A;
   input [23:0]B;
   output [47:0]Out;

   datapath i_0 (.B(B), .A(A), .Out(Out));
endmodule

module Reg(in, clk, out);
   input [31:0]in;
   input clk;
   output [31:0]out;

   DFF_X1 \out_reg[31]  (.D(in[31]), .CK(clk), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(in[30]), .CK(clk), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(in[29]), .CK(clk), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(in[28]), .CK(clk), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(in[27]), .CK(clk), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(in[26]), .CK(clk), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(in[25]), .CK(clk), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(in[24]), .CK(clk), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(in[23]), .CK(clk), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(in[22]), .CK(clk), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(in[21]), .CK(clk), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(in[20]), .CK(clk), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(in[19]), .CK(clk), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(in[18]), .CK(clk), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(in[17]), .CK(clk), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(in[16]), .CK(clk), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(in[15]), .CK(clk), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(in[14]), .CK(clk), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(in[13]), .CK(clk), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(in[12]), .CK(clk), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(in[11]), .CK(clk), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(in[10]), .CK(clk), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(in[9]), .CK(clk), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(in[8]), .CK(clk), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(in[7]), .CK(clk), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(in[6]), .CK(clk), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(in[5]), .CK(clk), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(in[4]), .CK(clk), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(in[3]), .CK(clk), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(in[2]), .CK(clk), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(in[1]), .CK(clk), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(in[0]), .CK(clk), .Q(out[0]), .QN());
endmodule

module datapath__0_4(p_0, p_1, MP_final);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]MP_final;

   XOR2_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .Z(MP_final[0]));
   AND2_X1 i_1 (.A1(p_1[0]), .A2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(p_1[1]), .B(n_0), .Z(MP_final[1]));
   AND2_X1 i_3 (.A1(n_0), .A2(p_1[1]), .ZN(n_1));
   XOR2_X1 i_4 (.A(p_1[2]), .B(n_1), .Z(MP_final[2]));
   AND2_X1 i_5 (.A1(n_1), .A2(p_1[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(p_1[3]), .B(n_2), .Z(MP_final[3]));
   AND2_X1 i_7 (.A1(n_2), .A2(p_1[3]), .ZN(n_3));
   XOR2_X1 i_8 (.A(p_1[4]), .B(n_3), .Z(MP_final[4]));
   AND2_X1 i_9 (.A1(n_3), .A2(p_1[4]), .ZN(n_4));
   XOR2_X1 i_10 (.A(p_1[5]), .B(n_4), .Z(MP_final[5]));
   AND2_X1 i_11 (.A1(n_4), .A2(p_1[5]), .ZN(n_5));
   XOR2_X1 i_12 (.A(p_1[6]), .B(n_5), .Z(MP_final[6]));
   AND2_X1 i_13 (.A1(n_5), .A2(p_1[6]), .ZN(n_6));
   XOR2_X1 i_14 (.A(p_1[7]), .B(n_6), .Z(MP_final[7]));
   AND2_X1 i_15 (.A1(n_6), .A2(p_1[7]), .ZN(n_7));
   XOR2_X1 i_16 (.A(p_1[8]), .B(n_7), .Z(MP_final[8]));
   AND2_X1 i_17 (.A1(n_7), .A2(p_1[8]), .ZN(n_8));
   XOR2_X1 i_18 (.A(p_1[9]), .B(n_8), .Z(MP_final[9]));
   AND2_X1 i_19 (.A1(n_8), .A2(p_1[9]), .ZN(n_9));
   XOR2_X1 i_20 (.A(p_1[10]), .B(n_9), .Z(MP_final[10]));
   AND2_X1 i_21 (.A1(n_9), .A2(p_1[10]), .ZN(n_10));
   XOR2_X1 i_22 (.A(p_1[11]), .B(n_10), .Z(MP_final[11]));
   AND2_X1 i_23 (.A1(n_10), .A2(p_1[11]), .ZN(n_11));
   XOR2_X1 i_24 (.A(p_1[12]), .B(n_11), .Z(MP_final[12]));
   AND2_X1 i_25 (.A1(n_11), .A2(p_1[12]), .ZN(n_12));
   XOR2_X1 i_26 (.A(p_1[13]), .B(n_12), .Z(MP_final[13]));
   XOR2_X1 i_28 (.A(p_1[14]), .B(n_21), .Z(MP_final[14]));
   XOR2_X1 i_30 (.A(p_1[15]), .B(n_20), .Z(MP_final[15]));
   XOR2_X1 i_32 (.A(p_1[16]), .B(n_19), .Z(MP_final[16]));
   XOR2_X1 i_34 (.A(p_1[17]), .B(n_18), .Z(MP_final[17]));
   XOR2_X1 i_36 (.A(p_1[18]), .B(n_17), .Z(MP_final[18]));
   XOR2_X1 i_38 (.A(p_1[19]), .B(n_16), .Z(MP_final[19]));
   XOR2_X1 i_40 (.A(p_1[20]), .B(n_15), .Z(MP_final[20]));
   XOR2_X1 i_42 (.A(p_1[21]), .B(n_14), .Z(MP_final[21]));
   XNOR2_X1 i_27 (.A(p_1[22]), .B(n_13), .ZN(MP_final[22]));
   NAND2_X1 i_29 (.A1(p_1[21]), .A2(n_14), .ZN(n_13));
   AND2_X1 i_31 (.A1(p_1[20]), .A2(n_15), .ZN(n_14));
   AND2_X1 i_33 (.A1(p_1[19]), .A2(n_16), .ZN(n_15));
   AND2_X1 i_35 (.A1(p_1[18]), .A2(n_17), .ZN(n_16));
   AND2_X1 i_37 (.A1(p_1[17]), .A2(n_18), .ZN(n_17));
   AND2_X1 i_39 (.A1(p_1[16]), .A2(n_19), .ZN(n_18));
   AND2_X1 i_41 (.A1(p_1[15]), .A2(n_20), .ZN(n_19));
   AND2_X1 i_43 (.A1(p_1[14]), .A2(n_21), .ZN(n_20));
   AND2_X1 i_44 (.A1(n_12), .A2(p_1[13]), .ZN(n_21));
endmodule

module float_mult(A, B, clk, Exception, Overflow, Underflow, Out);
   input [31:0]A;
   input [31:0]B;
   input clk;
   output Exception;
   output Overflow;
   output Underflow;
   output [31:0]Out;

   wire [31:0]afterB;
   wire [31:0]afterA;
   wire [47:0]MP;
   wire [22:0]MP_final;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_0_0;
   wire n_0_23;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_24;
   wire n_0_25;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_26;
   wire n_0_0_7;
   wire n_0_27;
   wire n_0_0_8;
   wire n_0_28;
   wire n_0_29;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_30;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_31;
   wire n_0_0_15;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_34;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_9;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_40;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_32;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_33;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_93;
   wire n_0_0_94;

   Reg__0_17 regB (.in(B), .clk(clk), .out(afterB));
   Reg__0_18 regA (.in(A), .clk(clk), .out(afterA));
   N_Bit_Mult mantissa_multiplier (.A({n_0_33, afterA[22], afterA[21], 
      afterA[20], afterA[19], afterA[18], afterA[17], afterA[16], afterA[15], 
      afterA[14], afterA[13], afterA[12], afterA[11], afterA[10], afterA[9], 
      afterA[8], afterA[7], afterA[6], afterA[5], afterA[4], afterA[3], 
      afterA[2], afterA[1], afterA[0]}), .B({n_0_32, afterB[22], afterB[21], 
      afterB[20], afterB[19], afterB[18], afterB[17], afterB[16], afterB[15], 
      afterB[14], afterB[13], afterB[12], afterB[11], afterB[10], afterB[9], 
      afterB[8], afterB[7], afterB[6], afterB[5], afterB[4], afterB[3], 
      afterB[2], afterB[1], afterB[0]}), .Out(MP));
   Reg regOut (.in({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0}), .clk(clk), .out(Out));
   datapath__0_4 i_0_6 (.p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, n_0_34}), .p_1({n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, 
      n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, 
      n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35}), 
      .MP_final(MP_final));
   AND2_X1 i_0_0_0 (.A1(MP_final[0]), .A2(n_0_0_0), .ZN(n_0_0));
   AND2_X1 i_0_0_1 (.A1(MP_final[1]), .A2(n_0_0_0), .ZN(n_0_1));
   AND2_X1 i_0_0_2 (.A1(MP_final[2]), .A2(n_0_0_0), .ZN(n_0_2));
   AND2_X1 i_0_0_3 (.A1(MP_final[3]), .A2(n_0_0_0), .ZN(n_0_3));
   AND2_X1 i_0_0_4 (.A1(MP_final[4]), .A2(n_0_0_0), .ZN(n_0_4));
   AND2_X1 i_0_0_5 (.A1(MP_final[5]), .A2(n_0_0_0), .ZN(n_0_5));
   AND2_X1 i_0_0_6 (.A1(MP_final[6]), .A2(n_0_0_0), .ZN(n_0_6));
   AND2_X1 i_0_0_7 (.A1(MP_final[7]), .A2(n_0_0_0), .ZN(n_0_7));
   AND2_X1 i_0_0_8 (.A1(MP_final[8]), .A2(n_0_0_0), .ZN(n_0_8));
   AND2_X1 i_0_0_9 (.A1(MP_final[9]), .A2(n_0_0_0), .ZN(n_0_9));
   AND2_X1 i_0_0_10 (.A1(MP_final[10]), .A2(n_0_0_0), .ZN(n_0_10));
   AND2_X1 i_0_0_11 (.A1(MP_final[11]), .A2(n_0_0_0), .ZN(n_0_11));
   AND2_X1 i_0_0_12 (.A1(MP_final[12]), .A2(n_0_0_0), .ZN(n_0_12));
   AND2_X1 i_0_0_13 (.A1(MP_final[13]), .A2(n_0_0_0), .ZN(n_0_13));
   AND2_X1 i_0_0_14 (.A1(MP_final[14]), .A2(n_0_0_0), .ZN(n_0_14));
   AND2_X1 i_0_0_15 (.A1(MP_final[15]), .A2(n_0_0_0), .ZN(n_0_15));
   AND2_X1 i_0_0_16 (.A1(MP_final[16]), .A2(n_0_0_0), .ZN(n_0_16));
   AND2_X1 i_0_0_17 (.A1(MP_final[17]), .A2(n_0_0_0), .ZN(n_0_17));
   AND2_X1 i_0_0_18 (.A1(MP_final[18]), .A2(n_0_0_0), .ZN(n_0_18));
   AND2_X1 i_0_0_19 (.A1(MP_final[19]), .A2(n_0_0_0), .ZN(n_0_19));
   AND2_X1 i_0_0_20 (.A1(MP_final[20]), .A2(n_0_0_0), .ZN(n_0_20));
   AND2_X1 i_0_0_21 (.A1(MP_final[21]), .A2(n_0_0_0), .ZN(n_0_21));
   AND2_X1 i_0_0_22 (.A1(MP_final[22]), .A2(n_0_0_0), .ZN(n_0_22));
   NOR2_X1 i_0_0_23 (.A1(n_0_0_39), .A2(n_0_0_12), .ZN(n_0_0_0));
   OAI21_X1 i_0_0_24 (.A(n_0_0_13), .B1(n_0_0_12), .B2(n_0_0_1), .ZN(n_0_23));
   XNOR2_X1 i_0_0_25 (.A(afterB[23]), .B(n_0_0_2), .ZN(n_0_0_1));
   XNOR2_X1 i_0_0_26 (.A(MP[47]), .B(afterA[23]), .ZN(n_0_0_2));
   OAI21_X1 i_0_0_27 (.A(n_0_0_13), .B1(n_0_0_12), .B2(n_0_0_18), .ZN(n_0_24));
   OAI21_X1 i_0_0_28 (.A(n_0_0_13), .B1(n_0_0_12), .B2(n_0_0_5), .ZN(n_0_25));
   XOR2_X1 i_0_0_29 (.A(n_0_0_54), .B(n_0_0_6), .Z(n_0_0_5));
   NAND2_X1 i_0_0_30 (.A1(n_0_0_53), .A2(n_0_0_55), .ZN(n_0_0_6));
   OAI33_X1 i_0_0_31 (.A1(Exception), .A2(n_0_0_35), .A3(n_0_0_26), .B1(n_0_0_12), 
      .B2(n_0_0_7), .B3(n_0_0_51), .ZN(n_0_26));
   AND2_X1 i_0_0_32 (.A1(n_0_0_58), .A2(n_0_0_52), .ZN(n_0_0_7));
   OAI21_X1 i_0_0_33 (.A(n_0_0_13), .B1(n_0_0_12), .B2(n_0_0_8), .ZN(n_0_27));
   XNOR2_X1 i_0_0_34 (.A(n_0_0_50), .B(n_0_0_47), .ZN(n_0_0_8));
   OAI21_X1 i_0_0_35 (.A(n_0_0_13), .B1(n_0_0_12), .B2(n_0_0_19), .ZN(n_0_28));
   OAI21_X1 i_0_0_36 (.A(n_0_0_13), .B1(n_0_0_12), .B2(n_0_0_10), .ZN(n_0_29));
   XNOR2_X1 i_0_0_37 (.A(n_0_0_45), .B(n_0_0_11), .ZN(n_0_0_10));
   AND2_X1 i_0_0_38 (.A1(n_0_0_72), .A2(n_0_0_71), .ZN(n_0_0_11));
   OAI21_X1 i_0_0_39 (.A(n_0_0_13), .B1(n_0_0_12), .B2(n_0_0_36), .ZN(n_0_30));
   OR2_X1 i_0_0_40 (.A1(n_0_0_38), .A2(n_0_0_14), .ZN(n_0_0_12));
   OR2_X1 i_0_0_41 (.A1(n_0_0_35), .A2(n_0_0_14), .ZN(n_0_0_13));
   OR2_X1 i_0_0_42 (.A1(n_0_0_26), .A2(Exception), .ZN(n_0_0_14));
   NOR2_X1 i_0_0_43 (.A1(Exception), .A2(n_0_0_15), .ZN(n_0_31));
   XNOR2_X1 i_0_0_44 (.A(afterB[31]), .B(afterA[31]), .ZN(n_0_0_15));
   NOR2_X1 i_0_0_45 (.A1(n_0_0_24), .A2(n_0_0_22), .ZN(Underflow));
   AOI21_X1 i_0_0_46 (.A(n_0_0_38), .B1(n_0_0_23), .B2(n_0_0_93), .ZN(n_0_0_22));
   NOR3_X1 i_0_0_47 (.A1(n_0_0_78), .A2(n_0_0_74), .A3(n_0_0_46), .ZN(n_0_0_23));
   NOR2_X1 i_0_0_48 (.A1(n_0_0_35), .A2(n_0_0_24), .ZN(Overflow));
   NOR2_X1 i_0_0_49 (.A1(Exception), .A2(n_0_0_25), .ZN(n_0_0_24));
   INV_X1 i_0_0_50 (.A(n_0_0_26), .ZN(n_0_0_25));
   NOR2_X1 i_0_0_51 (.A1(n_0_0_32), .A2(n_0_0_27), .ZN(n_0_0_26));
   NAND4_X1 i_0_0_52 (.A1(n_0_0_31), .A2(n_0_0_30), .A3(n_0_0_29), .A4(n_0_0_28), 
      .ZN(n_0_0_27));
   NOR4_X1 i_0_0_53 (.A1(MP_final[6]), .A2(MP_final[3]), .A3(MP_final[2]), 
      .A4(MP_final[0]), .ZN(n_0_0_28));
   NOR3_X1 i_0_0_54 (.A1(MP_final[5]), .A2(MP_final[4]), .A3(MP_final[1]), 
      .ZN(n_0_0_29));
   NOR4_X1 i_0_0_55 (.A1(MP_final[14]), .A2(MP_final[13]), .A3(MP_final[12]), 
      .A4(MP_final[11]), .ZN(n_0_0_30));
   NOR4_X1 i_0_0_56 (.A1(MP_final[10]), .A2(MP_final[9]), .A3(MP_final[8]), 
      .A4(MP_final[7]), .ZN(n_0_0_31));
   NAND2_X1 i_0_0_57 (.A1(n_0_0_34), .A2(n_0_0_33), .ZN(n_0_0_32));
   NOR4_X1 i_0_0_58 (.A1(MP_final[22]), .A2(MP_final[21]), .A3(MP_final[20]), 
      .A4(MP_final[19]), .ZN(n_0_0_33));
   NOR4_X1 i_0_0_59 (.A1(MP_final[18]), .A2(MP_final[17]), .A3(MP_final[16]), 
      .A4(MP_final[15]), .ZN(n_0_0_34));
   OAI21_X1 i_0_0_60 (.A(n_0_0_36), .B1(n_0_0_38), .B2(n_0_0_39), .ZN(n_0_0_35));
   XNOR2_X1 i_0_0_61 (.A(n_0_0_43), .B(n_0_0_37), .ZN(n_0_0_36));
   OR2_X1 i_0_0_62 (.A1(n_0_0_75), .A2(n_0_0_77), .ZN(n_0_0_37));
   NOR3_X1 i_0_0_63 (.A1(n_0_0_42), .A2(n_0_0_70), .A3(n_0_0_75), .ZN(n_0_0_38));
   NOR3_X1 i_0_0_64 (.A1(n_0_0_76), .A2(n_0_0_41), .A3(n_0_0_77), .ZN(n_0_0_39));
   NOR2_X1 i_0_0_65 (.A1(n_0_0_75), .A2(n_0_0_42), .ZN(n_0_0_41));
   INV_X1 i_0_0_66 (.A(n_0_0_43), .ZN(n_0_0_42));
   AND2_X1 i_0_0_67 (.A1(n_0_0_71), .A2(n_0_0_44), .ZN(n_0_0_43));
   NAND2_X1 i_0_0_68 (.A1(n_0_0_72), .A2(n_0_0_45), .ZN(n_0_0_44));
   OAI21_X1 i_0_0_69 (.A(n_0_0_46), .B1(n_0_0_21), .B2(n_0_0_49), .ZN(n_0_0_45));
   NAND2_X1 i_0_0_70 (.A1(n_0_0_40), .A2(n_0_0_20), .ZN(n_0_0_46));
   OR3_X1 i_0_0_71 (.A1(n_0_0_93), .A2(n_0_0_73), .A3(n_0_0_74), .ZN(n_0_0_71));
   OAI21_X1 i_0_0_72 (.A(n_0_0_74), .B1(n_0_0_73), .B2(n_0_0_93), .ZN(n_0_0_72));
   NOR2_X1 i_0_0_73 (.A1(afterB[29]), .A2(afterA[29]), .ZN(n_0_0_73));
   NAND2_X1 i_0_0_74 (.A1(afterB[28]), .A2(afterA[28]), .ZN(n_0_0_74));
   AOI21_X1 i_0_0_75 (.A(n_0_0_94), .B1(n_0_0_70), .B2(n_0_0_78), .ZN(n_0_0_75));
   OAI21_X1 i_0_0_76 (.A(n_0_0_80), .B1(n_0_0_79), .B2(MP[47]), .ZN(n_0_34));
   NAND2_X1 i_0_0_77 (.A1(n_0_0_81), .A2(MP[22]), .ZN(n_0_0_79));
   OAI211_X1 i_0_0_78 (.A(MP[47]), .B(MP[23]), .C1(n_0_0_81), .C2(MP[22]), 
      .ZN(n_0_0_80));
   NAND3_X1 i_0_0_79 (.A1(n_0_0_88), .A2(n_0_0_87), .A3(n_0_0_82), .ZN(n_0_0_81));
   AND4_X1 i_0_0_80 (.A1(n_0_0_86), .A2(n_0_0_85), .A3(n_0_0_84), .A4(n_0_0_83), 
      .ZN(n_0_0_82));
   NOR4_X1 i_0_0_81 (.A1(MP[7]), .A2(MP[6]), .A3(MP[5]), .A4(MP[4]), .ZN(
      n_0_0_83));
   NOR4_X1 i_0_0_82 (.A1(MP[3]), .A2(MP[2]), .A3(MP[1]), .A4(MP[0]), .ZN(
      n_0_0_84));
   NOR4_X1 i_0_0_83 (.A1(MP[15]), .A2(MP[14]), .A3(MP[13]), .A4(MP[12]), 
      .ZN(n_0_0_85));
   NOR4_X1 i_0_0_84 (.A1(MP[11]), .A2(MP[10]), .A3(MP[9]), .A4(MP[8]), .ZN(
      n_0_0_86));
   NOR4_X1 i_0_0_85 (.A1(MP[19]), .A2(MP[18]), .A3(MP[17]), .A4(MP[16]), 
      .ZN(n_0_0_87));
   NOR2_X1 i_0_0_86 (.A1(MP[21]), .A2(MP[20]), .ZN(n_0_0_88));
   MUX2_X1 i_0_0_126 (.A(MP[23]), .B(MP[24]), .S(MP[47]), .Z(n_0_35));
   MUX2_X1 i_0_0_127 (.A(MP[24]), .B(MP[25]), .S(MP[47]), .Z(n_0_36));
   MUX2_X1 i_0_0_128 (.A(MP[25]), .B(MP[26]), .S(MP[47]), .Z(n_0_37));
   MUX2_X1 i_0_0_129 (.A(MP[26]), .B(MP[27]), .S(MP[47]), .Z(n_0_38));
   MUX2_X1 i_0_0_130 (.A(MP[27]), .B(MP[28]), .S(MP[47]), .Z(n_0_39));
   MUX2_X1 i_0_0_131 (.A(MP[28]), .B(MP[29]), .S(MP[47]), .Z(n_0_40));
   MUX2_X1 i_0_0_132 (.A(MP[29]), .B(MP[30]), .S(MP[47]), .Z(n_0_41));
   MUX2_X1 i_0_0_133 (.A(MP[30]), .B(MP[31]), .S(MP[47]), .Z(n_0_42));
   MUX2_X1 i_0_0_134 (.A(MP[31]), .B(MP[32]), .S(MP[47]), .Z(n_0_43));
   MUX2_X1 i_0_0_135 (.A(MP[32]), .B(MP[33]), .S(MP[47]), .Z(n_0_44));
   MUX2_X1 i_0_0_136 (.A(MP[33]), .B(MP[34]), .S(MP[47]), .Z(n_0_45));
   MUX2_X1 i_0_0_137 (.A(MP[34]), .B(MP[35]), .S(MP[47]), .Z(n_0_46));
   MUX2_X1 i_0_0_138 (.A(MP[35]), .B(MP[36]), .S(MP[47]), .Z(n_0_47));
   MUX2_X1 i_0_0_139 (.A(MP[36]), .B(MP[37]), .S(MP[47]), .Z(n_0_48));
   MUX2_X1 i_0_0_140 (.A(MP[37]), .B(MP[38]), .S(MP[47]), .Z(n_0_49));
   MUX2_X1 i_0_0_141 (.A(MP[38]), .B(MP[39]), .S(MP[47]), .Z(n_0_50));
   MUX2_X1 i_0_0_142 (.A(MP[39]), .B(MP[40]), .S(MP[47]), .Z(n_0_51));
   MUX2_X1 i_0_0_143 (.A(MP[40]), .B(MP[41]), .S(MP[47]), .Z(n_0_52));
   MUX2_X1 i_0_0_144 (.A(MP[41]), .B(MP[42]), .S(MP[47]), .Z(n_0_53));
   MUX2_X1 i_0_0_145 (.A(MP[42]), .B(MP[43]), .S(MP[47]), .Z(n_0_54));
   MUX2_X1 i_0_0_146 (.A(MP[43]), .B(MP[44]), .S(MP[47]), .Z(n_0_55));
   MUX2_X1 i_0_0_147 (.A(MP[44]), .B(MP[45]), .S(MP[47]), .Z(n_0_56));
   MUX2_X1 i_0_0_148 (.A(MP[45]), .B(MP[46]), .S(MP[47]), .Z(n_0_57));
   OAI22_X1 i_0_0_87 (.A1(n_0_0_92), .A2(n_0_0_91), .B1(n_0_0_90), .B2(n_0_0_89), 
      .ZN(Exception));
   NAND4_X1 i_0_0_88 (.A1(afterA[30]), .A2(afterA[29]), .A3(afterA[28]), 
      .A4(afterA[27]), .ZN(n_0_0_89));
   NAND4_X1 i_0_0_89 (.A1(afterA[26]), .A2(afterA[25]), .A3(afterA[24]), 
      .A4(afterA[23]), .ZN(n_0_0_90));
   NAND4_X1 i_0_0_90 (.A1(afterB[30]), .A2(afterB[29]), .A3(afterB[28]), 
      .A4(afterB[27]), .ZN(n_0_0_91));
   NAND4_X1 i_0_0_91 (.A1(afterB[26]), .A2(afterB[25]), .A3(afterB[24]), 
      .A4(afterB[23]), .ZN(n_0_0_92));
   NAND3_X1 i_0_0_92 (.A1(afterB[23]), .A2(MP[47]), .A3(afterA[23]), .ZN(n_0_0_3));
   NOR3_X1 i_0_0_93 (.A1(afterB[23]), .A2(MP[47]), .A3(afterA[23]), .ZN(n_0_0_4));
   XNOR2_X1 i_0_0_94 (.A(afterB[24]), .B(afterA[24]), .ZN(n_0_0_9));
   INV_X1 i_0_0_95 (.A(n_0_0_4), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_96 (.A1(n_0_0_16), .A2(n_0_0_3), .ZN(n_0_0_17));
   XNOR2_X1 i_0_0_97 (.A(n_0_0_9), .B(n_0_0_17), .ZN(n_0_0_18));
   XNOR2_X1 i_0_0_98 (.A(n_0_0_40), .B(n_0_0_20), .ZN(n_0_0_19));
   XOR2_X1 i_0_0_99 (.A(n_0_0_49), .B(n_0_0_21), .Z(n_0_0_20));
   XNOR2_X1 i_0_0_100 (.A(afterB[28]), .B(afterA[28]), .ZN(n_0_0_21));
   OAI22_X1 i_0_0_101 (.A1(n_0_0_62), .A2(n_0_0_48), .B1(n_0_0_50), .B2(n_0_0_47), 
      .ZN(n_0_0_40));
   XNOR2_X1 i_0_0_102 (.A(n_0_0_62), .B(n_0_0_48), .ZN(n_0_0_47));
   OAI21_X1 i_0_0_103 (.A(n_0_0_49), .B1(afterB[27]), .B2(afterA[27]), .ZN(
      n_0_0_48));
   NAND2_X1 i_0_0_104 (.A1(afterB[27]), .A2(afterA[27]), .ZN(n_0_0_49));
   NOR2_X1 i_0_0_105 (.A1(n_0_0_60), .A2(n_0_0_51), .ZN(n_0_0_50));
   NOR2_X1 i_0_0_106 (.A1(n_0_0_58), .A2(n_0_0_52), .ZN(n_0_0_51));
   AOI21_X1 i_0_0_107 (.A(n_0_0_56), .B1(n_0_0_54), .B2(n_0_0_53), .ZN(n_0_0_52));
   OAI21_X1 i_0_0_108 (.A(n_0_0_57), .B1(n_0_0_65), .B2(n_0_0_64), .ZN(n_0_0_53));
   AOI21_X1 i_0_0_109 (.A(n_0_0_4), .B1(n_0_0_9), .B2(n_0_0_3), .ZN(n_0_0_54));
   INV_X1 i_0_0_110 (.A(n_0_0_56), .ZN(n_0_0_55));
   NOR3_X1 i_0_0_111 (.A1(n_0_0_65), .A2(n_0_0_64), .A3(n_0_0_57), .ZN(n_0_0_56));
   OAI21_X1 i_0_0_112 (.A(n_0_0_63), .B1(afterB[25]), .B2(afterA[25]), .ZN(
      n_0_0_57));
   INV_X1 i_0_0_113 (.A(n_0_0_59), .ZN(n_0_0_58));
   AOI21_X1 i_0_0_114 (.A(n_0_0_60), .B1(n_0_0_63), .B2(n_0_0_61), .ZN(n_0_0_59));
   NOR2_X1 i_0_0_115 (.A1(n_0_0_63), .A2(n_0_0_61), .ZN(n_0_0_60));
   OAI21_X1 i_0_0_116 (.A(n_0_0_62), .B1(afterB[26]), .B2(afterA[26]), .ZN(
      n_0_0_61));
   NAND2_X1 i_0_0_117 (.A1(afterB[26]), .A2(afterA[26]), .ZN(n_0_0_62));
   NAND2_X1 i_0_0_118 (.A1(afterB[25]), .A2(afterA[25]), .ZN(n_0_0_63));
   INV_X1 i_0_0_119 (.A(afterA[24]), .ZN(n_0_0_64));
   INV_X1 i_0_0_120 (.A(afterB[24]), .ZN(n_0_0_65));
   NAND2_X1 i_0_0_121 (.A1(n_0_0_67), .A2(n_0_0_66), .ZN(n_0_32));
   NOR4_X1 i_0_0_122 (.A1(afterB[25]), .A2(afterB[24]), .A3(afterB[30]), 
      .A4(afterB[27]), .ZN(n_0_0_66));
   NOR4_X1 i_0_0_123 (.A1(afterB[26]), .A2(afterB[23]), .A3(afterB[29]), 
      .A4(afterB[28]), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_124 (.A1(n_0_0_69), .A2(n_0_0_68), .ZN(n_0_33));
   NOR4_X1 i_0_0_125 (.A1(afterA[25]), .A2(afterA[24]), .A3(afterA[30]), 
      .A4(afterA[27]), .ZN(n_0_0_68));
   NOR4_X1 i_0_0_149 (.A1(afterA[26]), .A2(afterA[23]), .A3(afterA[29]), 
      .A4(afterA[28]), .ZN(n_0_0_69));
   INV_X1 i_0_0_150 (.A(n_0_0_76), .ZN(n_0_0_70));
   NOR2_X1 i_0_0_151 (.A1(afterB[30]), .A2(afterA[30]), .ZN(n_0_0_76));
   AND3_X1 i_0_0_152 (.A1(n_0_0_70), .A2(n_0_0_78), .A3(n_0_0_94), .ZN(n_0_0_77));
   NAND2_X1 i_0_0_153 (.A1(afterB[30]), .A2(afterA[30]), .ZN(n_0_0_78));
   INV_X1 i_0_0_154 (.A(n_0_0_94), .ZN(n_0_0_93));
   NAND2_X1 i_0_0_155 (.A1(afterB[29]), .A2(afterA[29]), .ZN(n_0_0_94));
endmodule
