/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Jan  4 05:03:18 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3461303721 */

module datapath(p_0, p_1);
   output [63:0]p_0;
   input [63:0]p_1;

   XOR2_X1 i_0 (.A(p_1[1]), .B(p_1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(p_1[2]), .B1(p_1[1]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(p_1[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(p_1[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(p_1[6]), .B1(n_27), .B2(p_1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(p_1[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(p_1[9]), .B1(n_25), .B2(p_1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(p_1[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(p_1[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(p_1[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(p_1[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(p_1[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(p_1[16]), .B1(n_19), .B2(p_1[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(p_1[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(p_1[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(p_1[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(p_1[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(p_1[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(p_1[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(p_1[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(p_1[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(p_1[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(p_1[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(p_1[27]), .B1(n_9), .B2(p_1[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(p_1[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(p_1[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(p_1[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(p_1[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .A4(p_1[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(p_1[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(p_1[26]), .A3(p_1[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(p_1[23]), .A3(p_1[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(p_1[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(p_1[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .A4(p_1[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(p_1[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(p_1[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(p_1[15]), .A3(p_1[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(p_1[12]), .A3(p_1[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(p_1[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(p_1[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(p_1[8]), .A3(p_1[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(p_1[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(p_1[5]), .A3(p_1[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(p_1[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(p_1[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(p_1[2]), .A2(p_1[1]), .A3(p_1[0]), .ZN(n_29));
   INV_X1 i_61 (.A(p_1[11]), .ZN(n_30));
   INV_X1 i_62 (.A(p_1[14]), .ZN(n_31));
   INV_X1 i_63 (.A(p_1[21]), .ZN(n_32));
   INV_X1 i_64 (.A(p_1[25]), .ZN(n_33));
endmodule

module halfadder__1_1873(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1874(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_1873 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_1865(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1862(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1866(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1865 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1862 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1857(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1854(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1858(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1857 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1854 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1849(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1846(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1850(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1849 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1846 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1841(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1838(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1842(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1841 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1838 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1833(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1830(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1833 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1830 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1825(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1822(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1826(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1825 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1822 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1817(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1814(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1817 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1814 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1809(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1806(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1809 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1806 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1801(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1798(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1802(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1801 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1798 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1793(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1790(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1793 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1790 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1782(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1785 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1782 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1778(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1777 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1774 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1769 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1766 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1761 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1758 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1750(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1753 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1750 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1745(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1742(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1745 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1742 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1737(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1734(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1737 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1734 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1729(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1726(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1730(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1729 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1726 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1721(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1718(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1722(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1721 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1718 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1713(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1710(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1714(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1713 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1710 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1705(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1702(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1706(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1705 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1702 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1697(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1694(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1698(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1697 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1694 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1689(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1686(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1690(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1689 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1686 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1681(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1678(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1682(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1681 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1678 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1673(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1670(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1674(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1673 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1670 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1665(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1662(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1666(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1665 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1662 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1657(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1654(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1658(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1657 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1654 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1649(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1646(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1650(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1649 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1646 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1641(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1638(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1642(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1641 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1638 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1633(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1630(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1634(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1633 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1630 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1625(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1622(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1626(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1625 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1622 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1617(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1614(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1618(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1617 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1614 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1609(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1606(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1610(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1609 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1606 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1601(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1598(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1602(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1601 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1598 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1593(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1590(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1594(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1593 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1590 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1585(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1582(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1586(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1585 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1582 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1577(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1574(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1578(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1577 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1574 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1569(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1566(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1570(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1569 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1566 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1561(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1558(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1562(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1561 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1558 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1553(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1550(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1554(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1553 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1550 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1545(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1542(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1546(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1545 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1542 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1537(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1534(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1538(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1537 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1534 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1530(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1529 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1526 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_1518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_1522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_1521 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_1518 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__1_1369(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1370(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_1369 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_1361(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1358(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1362(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1361 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1358 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1353(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1350(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1354(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1353 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1350 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1345(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1342(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1346(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1345 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1342 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1337(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1334(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1337 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1334 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1329(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1326(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1330(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1329 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1326 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1321(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1318(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1322(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1321 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1318 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1313(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1310(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1313 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1310 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1305(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1302(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1306(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1305 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1302 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1297(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1294(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1298(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1297 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1294 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1289(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1286(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1289 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1286 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1278(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1281 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1278 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1273 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1270 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1265 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1262 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1258(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1257 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1254 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1246(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1249 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1246 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1241(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1238(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1241 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1238 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1233(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1230(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1234(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1233 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1230 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1225(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1222(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1226(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1225 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1222 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1217(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1214(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1217 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1214 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1209(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1206(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1210(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1209 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1206 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1201(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1198(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1202(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1201 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1198 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1193(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1190(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1194(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1193 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1190 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1185(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1182(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1186(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1185 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1182 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1177(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1174(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1178(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1177 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1174 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1169(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1166(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1170(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1169 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1166 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1161(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1158(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1162(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1161 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1158 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1153(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1150(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1154(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1153 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1150 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1145(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1142(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1146(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1145 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1142 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1137(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1134(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1138(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1137 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1134 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1129(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1126(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1130(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1129 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1126 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1121(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1118(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1122(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1121 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1118 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1113(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1110(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1114(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1113 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1110 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1105(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1102(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1106(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1105 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1102 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1097(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1094(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1098(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1097 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1094 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1089(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1086(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1090(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1089 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1086 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1081(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1078(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1082(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1081 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1078 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1073(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1070(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1074(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1073 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1070 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1065(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1062(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1066(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1065 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1062 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1057(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1054(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1058(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1057 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1054 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1049(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1046(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1050(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1049 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1046 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1041(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1038(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1042(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1041 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1038 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1033(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1030(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1034(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1033 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1030 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1025(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_1022(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_1026(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_1025 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_1022 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__1_2043(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__1_1874 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(), .sum(s[19]), 
      .carry(c1[19]));
   fulladder__1_1866 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(
      s1[20]), .carry(c1[20]));
   fulladder__1_1858 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(
      s1[21]), .carry(c1[21]));
   fulladder__1_1850 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(
      s1[22]), .carry(c1[22]));
   fulladder__1_1842 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__1_1834 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__1_1826 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__1_1818 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__1_1810 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__1_1802 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__1_1794 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__1_1786 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__1_1778 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__1_1770 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__1_1762 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__1_1754 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__1_1746 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__1_1738 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__1_1730 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__1_1722 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__1_1714 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__1_1706 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__1_1698 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__1_1690 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__1_1682 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__1_1674 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__1_1666 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__1_1658 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__1_1650 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__1_1642 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__1_1634 genblk1_49_a (.a(x[63]), .b(y[49]), .cin(z[49]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__1_1626 genblk1_50_a (.a(x[63]), .b(y[63]), .cin(z[50]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__1_1618 genblk1_51_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__1_1610 genblk1_52_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__1_1602 genblk1_53_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__1_1594 genblk1_54_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__1_1586 genblk1_55_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__1_1578 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__1_1570 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__1_1562 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__1_1554 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__1_1546 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__1_1538 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__1_1530 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__1_1522 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__1_1370 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(), .sum(s[20]), 
      .carry(c2[20]));
   fulladder__1_1362 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), 
      .sum(s[21]), .carry(c2[21]));
   fulladder__1_1354 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), 
      .sum(s[22]), .carry(c2[22]));
   fulladder__1_1346 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), 
      .sum(s[23]), .carry(c2[23]));
   fulladder__1_1338 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__1_1330 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__1_1322 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__1_1314 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__1_1306 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__1_1298 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__1_1290 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__1_1282 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__1_1274 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__1_1266 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__1_1258 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__1_1250 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__1_1242 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__1_1234 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__1_1226 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__1_1218 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__1_1210 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__1_1202 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__1_1194 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__1_1186 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__1_1178 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__1_1170 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__1_1162 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__1_1154 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__1_1146 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__1_1138 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__1_1130 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__1_1122 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__1_1114 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__1_1106 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__1_1098 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__1_1090 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__1_1082 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__1_1074 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__1_1066 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__1_1058 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__1_1050 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__1_1042 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__1_1034 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__1_1026 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__1_3042(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3043(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_3042 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_3034(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3031(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3035(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3034 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3031 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3026(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3023(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3027(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3026 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3023 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3018(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3015(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3019(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3018 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3015 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3010(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3007(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3011(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3010 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3007 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3002(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2999(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3003(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3002 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2999 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2994(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2991(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2995(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2994 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2991 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2986(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2983(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2987(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2986 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2983 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2978(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2975(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2979(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2978 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2975 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2970(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2967(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2971(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2970 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2967 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2962(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2959(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2963(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2962 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2959 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2954(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2951(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2955(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2954 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2951 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2946(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2943(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2947(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2946 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2943 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2938(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2935(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2939(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2938 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2935 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2930(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2927(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2931(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2930 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2927 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2922(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2919(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2923(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2922 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2919 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2914(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2911(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2915(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2914 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2911 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2906(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2903(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2907(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2906 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2903 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2898(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2895(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2899(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2898 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2895 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2890(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2887(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2891(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2890 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2887 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2882(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2879(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2883(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2882 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2879 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2874(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2871(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2875(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2874 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2871 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2866(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2863(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2867(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2866 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2863 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2858(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2855(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2859(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2858 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2855 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2850(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2847(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2851(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2850 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2847 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2842(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2839(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2843(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2842 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2839 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2834(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2831(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2835(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2834 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2831 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2826(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2823(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2827(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2826 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2823 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2818(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2815(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2819(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2818 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2815 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2810(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2807(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2811(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2810 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2807 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2802(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2799(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2803(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2802 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2799 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2794(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2791(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2795(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2794 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2791 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2786(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2783(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2787(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2786 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2783 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2778(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2775(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2779(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2778 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2775 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2770(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2767(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2771(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2770 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2767 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2762(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2759(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2763(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2762 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2759 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2754(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2751(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2755(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2754 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2751 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2746(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2743(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2747(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2746 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2743 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2738(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2735(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2739(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2738 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2735 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2730(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2727(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2731(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2730 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2727 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2722(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2719(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2723(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2722 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2719 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2714(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2711(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2715(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2714 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2711 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2706(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2703(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2707(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2706 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2703 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2698(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2695(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2699(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2698 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2695 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2690(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2687(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2691(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2690 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2687 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2682(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2679(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2683(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2682 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2679 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2674(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2671(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2675(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2674 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2671 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2666(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2663(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2667(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2666 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2663 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2658(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2655(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2659(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2658 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2655 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2650(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2647(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2651(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2650 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2647 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2642(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2639(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2643(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2642 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2639 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2634(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2631(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2635(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2634 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2631 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2626(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2623(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2627(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2626 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2623 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2618(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2615(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2619(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2618 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2615 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2610(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2607(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2611(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2610 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2607 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2602(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2599(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2603(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2602 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2599 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2594(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2591(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2595(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2594 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2591 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2586(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2583(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2587(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2586 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2583 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2578(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2575(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2579(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2578 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2575 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2570(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2567(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2571(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2570 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2567 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2562(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2559(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2563(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2562 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2559 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2554(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2551(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2555(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2554 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2551 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2546(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_2543(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_2547(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_2546 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_2543 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__1_2538(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2539(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_2538 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_2530(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2527(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2531(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2530 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2527 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2522(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2519(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2523(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2522 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2519 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2514(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2511(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2515(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2514 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2511 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2506(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2503(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2507(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2506 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2503 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2498(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2495(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2499(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2498 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2495 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2490(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2487(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2491(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2490 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2487 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2482(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2479(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2483(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2482 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2479 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2474(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2471(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2475(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2474 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2471 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2466(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2463(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2467(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2466 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2463 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2458(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2455(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2459(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2458 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2455 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2450(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2447(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2451(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2450 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2447 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2442(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2439(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2443(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2442 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2439 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2434(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2431(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2435(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2434 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2431 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2426(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2423(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2427(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2426 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2423 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2418(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2415(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2419(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2418 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2415 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2410(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2407(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2411(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2410 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2407 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2402(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2399(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2403(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2402 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2399 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2394(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2391(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2395(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2394 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2391 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2386(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2383(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2387(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2386 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2383 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2378(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2375(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2379(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2378 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2375 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2370(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2367(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2371(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2370 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2367 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2362(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2359(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2363(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2362 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2359 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2354(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2351(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2355(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2354 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2351 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2346(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2343(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2347(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2346 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2343 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2338(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2335(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2339(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2338 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2335 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2330(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2327(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2331(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2330 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2327 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2322(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2319(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2323(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2322 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2319 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2314(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2311(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2315(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2314 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2311 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2306(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2303(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2307(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2306 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2303 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2298(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2295(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2299(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2298 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2295 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2290(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2287(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2291(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2290 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2287 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2282(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2279(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2283(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2282 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2279 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2274(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2271(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2275(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2274 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2271 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2266(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2263(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2267(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2266 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2263 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2258(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2255(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2259(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2258 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2255 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2250(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2247(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2251(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2250 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2247 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2242(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2239(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2243(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2242 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2239 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2234(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2231(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2235(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2234 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2231 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2226(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2223(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2227(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2226 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2223 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2218(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2215(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2219(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2218 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2215 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2210(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2207(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2211(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2210 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2207 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2202(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2199(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2203(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2202 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2199 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2194(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2191(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2195(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2194 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2191 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2186(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2183(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2187(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2186 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2183 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2178(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2175(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2179(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2178 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2175 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2170(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2167(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2171(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2170 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2167 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2162(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2159(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2163(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2162 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2159 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2154(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2151(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2155(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2154 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2151 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2146(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2143(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2147(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2146 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2143 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2138(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2135(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2139(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2138 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2135 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2130(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2127(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2131(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2130 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2127 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2122(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2119(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2123(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2122 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2119 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2114(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2111(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2115(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2114 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2111 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2106(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2103(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2107(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2106 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2103 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2098(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2095(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2099(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2098 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2095 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2090(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2087(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2091(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2090 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2087 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2082(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2079(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2083(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2082 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2079 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2074(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2071(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2075(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2074 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2071 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2066(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2063(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2067(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2066 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2063 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2058(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_2055(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_2059(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_2058 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_2055 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2050(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_2047(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_2051(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_2050 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_2047 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__1_3068(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__1_3043 genblk1_1_a (.a(x[1]), .b(y[1]), .cin(), .sum(s[1]), 
      .carry(c1[1]));
   fulladder__1_3035 genblk1_2_a (.a(x[2]), .b(y[2]), .cin(z[2]), .sum(s1[2]), 
      .carry(c1[2]));
   fulladder__1_3027 genblk1_3_a (.a(x[3]), .b(y[3]), .cin(z[3]), .sum(s1[3]), 
      .carry(c1[3]));
   fulladder__1_3019 genblk1_4_a (.a(x[4]), .b(y[4]), .cin(z[4]), .sum(s1[4]), 
      .carry(c1[4]));
   fulladder__1_3011 genblk1_5_a (.a(x[5]), .b(y[5]), .cin(z[5]), .sum(s1[5]), 
      .carry(c1[5]));
   fulladder__1_3003 genblk1_6_a (.a(x[6]), .b(y[6]), .cin(z[6]), .sum(s1[6]), 
      .carry(c1[6]));
   fulladder__1_2995 genblk1_7_a (.a(x[7]), .b(y[7]), .cin(z[7]), .sum(s1[7]), 
      .carry(c1[7]));
   fulladder__1_2987 genblk1_8_a (.a(x[8]), .b(y[8]), .cin(z[8]), .sum(s1[8]), 
      .carry(c1[8]));
   fulladder__1_2979 genblk1_9_a (.a(x[9]), .b(y[9]), .cin(z[9]), .sum(s1[9]), 
      .carry(c1[9]));
   fulladder__1_2971 genblk1_10_a (.a(x[10]), .b(y[10]), .cin(z[10]), .sum(
      s1[10]), .carry(c1[10]));
   fulladder__1_2963 genblk1_11_a (.a(x[11]), .b(y[11]), .cin(z[11]), .sum(
      s1[11]), .carry(c1[11]));
   fulladder__1_2955 genblk1_12_a (.a(x[12]), .b(y[12]), .cin(z[12]), .sum(
      s1[12]), .carry(c1[12]));
   fulladder__1_2947 genblk1_13_a (.a(x[13]), .b(y[13]), .cin(z[13]), .sum(
      s1[13]), .carry(c1[13]));
   fulladder__1_2939 genblk1_14_a (.a(x[14]), .b(y[14]), .cin(z[14]), .sum(
      s1[14]), .carry(c1[14]));
   fulladder__1_2931 genblk1_15_a (.a(x[15]), .b(y[15]), .cin(z[15]), .sum(
      s1[15]), .carry(c1[15]));
   fulladder__1_2923 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(z[16]), .sum(
      s1[16]), .carry(c1[16]));
   fulladder__1_2915 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(z[17]), .sum(
      s1[17]), .carry(c1[17]));
   fulladder__1_2907 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(
      s1[18]), .carry(c1[18]));
   fulladder__1_2899 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(
      s1[19]), .carry(c1[19]));
   fulladder__1_2891 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(
      s1[20]), .carry(c1[20]));
   fulladder__1_2883 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(
      s1[21]), .carry(c1[21]));
   fulladder__1_2875 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(
      s1[22]), .carry(c1[22]));
   fulladder__1_2867 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__1_2859 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__1_2851 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__1_2843 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__1_2835 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__1_2827 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__1_2819 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__1_2811 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__1_2803 genblk1_31_a (.a(x[63]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__1_2795 genblk1_32_a (.a(x[63]), .b(y[63]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__1_2787 genblk1_33_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__1_2779 genblk1_34_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__1_2771 genblk1_35_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__1_2763 genblk1_36_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__1_2755 genblk1_37_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__1_2747 genblk1_38_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__1_2739 genblk1_39_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__1_2731 genblk1_40_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__1_2723 genblk1_41_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__1_2715 genblk1_42_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__1_2707 genblk1_43_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__1_2699 genblk1_44_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__1_2691 genblk1_45_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__1_2683 genblk1_46_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__1_2675 genblk1_47_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__1_2667 genblk1_48_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__1_2659 genblk1_49_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__1_2651 genblk1_50_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__1_2643 genblk1_51_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__1_2635 genblk1_52_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__1_2627 genblk1_53_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__1_2619 genblk1_54_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__1_2611 genblk1_55_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__1_2603 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__1_2595 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__1_2587 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__1_2579 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__1_2571 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__1_2563 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__1_2555 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__1_2547 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__1_2539 genblk2_1_b (.a(s1[2]), .b(c1[1]), .cin(), .sum(s[2]), 
      .carry(c2[2]));
   fulladder__1_2531 genblk2_2_b (.a(s1[3]), .b(c1[2]), .cin(c2[2]), .sum(s[3]), 
      .carry(c2[3]));
   fulladder__1_2523 genblk2_3_b (.a(s1[4]), .b(c1[3]), .cin(c2[3]), .sum(s[4]), 
      .carry(c2[4]));
   fulladder__1_2515 genblk2_4_b (.a(s1[5]), .b(c1[4]), .cin(c2[4]), .sum(s[5]), 
      .carry(c2[5]));
   fulladder__1_2507 genblk2_5_b (.a(s1[6]), .b(c1[5]), .cin(c2[5]), .sum(s[6]), 
      .carry(c2[6]));
   fulladder__1_2499 genblk2_6_b (.a(s1[7]), .b(c1[6]), .cin(c2[6]), .sum(s[7]), 
      .carry(c2[7]));
   fulladder__1_2491 genblk2_7_b (.a(s1[8]), .b(c1[7]), .cin(c2[7]), .sum(s[8]), 
      .carry(c2[8]));
   fulladder__1_2483 genblk2_8_b (.a(s1[9]), .b(c1[8]), .cin(c2[8]), .sum(s[9]), 
      .carry(c2[9]));
   fulladder__1_2475 genblk2_9_b (.a(s1[10]), .b(c1[9]), .cin(c2[9]), .sum(s[10]), 
      .carry(c2[10]));
   fulladder__1_2467 genblk2_10_b (.a(s1[11]), .b(c1[10]), .cin(c2[10]), 
      .sum(s[11]), .carry(c2[11]));
   fulladder__1_2459 genblk2_11_b (.a(s1[12]), .b(c1[11]), .cin(c2[11]), 
      .sum(s[12]), .carry(c2[12]));
   fulladder__1_2451 genblk2_12_b (.a(s1[13]), .b(c1[12]), .cin(c2[12]), 
      .sum(s[13]), .carry(c2[13]));
   fulladder__1_2443 genblk2_13_b (.a(s1[14]), .b(c1[13]), .cin(c2[13]), 
      .sum(s[14]), .carry(c2[14]));
   fulladder__1_2435 genblk2_14_b (.a(s1[15]), .b(c1[14]), .cin(c2[14]), 
      .sum(s[15]), .carry(c2[15]));
   fulladder__1_2427 genblk2_15_b (.a(s1[16]), .b(c1[15]), .cin(c2[15]), 
      .sum(s[16]), .carry(c2[16]));
   fulladder__1_2419 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(c2[16]), 
      .sum(s[17]), .carry(c2[17]));
   fulladder__1_2411 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), 
      .sum(s[18]), .carry(c2[18]));
   fulladder__1_2403 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), 
      .sum(s[19]), .carry(c2[19]));
   fulladder__1_2395 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), 
      .sum(s[20]), .carry(c2[20]));
   fulladder__1_2387 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), 
      .sum(s[21]), .carry(c2[21]));
   fulladder__1_2379 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), 
      .sum(s[22]), .carry(c2[22]));
   fulladder__1_2371 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), 
      .sum(s[23]), .carry(c2[23]));
   fulladder__1_2363 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__1_2355 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__1_2347 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__1_2339 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__1_2331 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__1_2323 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__1_2315 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__1_2307 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__1_2299 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__1_2291 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__1_2283 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__1_2275 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__1_2267 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__1_2259 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__1_2251 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__1_2243 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__1_2235 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__1_2227 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__1_2219 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__1_2211 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__1_2203 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__1_2195 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__1_2187 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__1_2179 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__1_2171 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__1_2163 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__1_2155 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__1_2147 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__1_2139 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__1_2131 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__1_2123 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__1_2115 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__1_2107 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__1_2099 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__1_2091 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__1_2083 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__1_2075 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__1_2067 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__1_2059 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__1_2051 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__1_4043(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4044(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_4043 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_4035(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4032(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4036(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4035 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4032 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4027(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4024(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4028(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4027 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4024 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4019(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4016(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4020(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4019 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4016 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4011(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4008(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4012(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4011 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4008 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4003(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4000(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4004(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4003 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4000 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3995(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3992(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3996(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3995 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3992 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3987(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3984(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3988(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3987 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3984 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3979(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3976(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3980(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3979 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3976 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3971(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3968(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3972(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3971 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3968 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3963(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3960(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3964(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3963 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3960 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3955(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3952(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3956(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3955 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3952 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3947(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3944(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3948(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3947 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3944 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3939(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3936(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3940(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3939 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3936 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3931(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3928(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3932(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3931 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3928 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3923(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3920(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3924(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3923 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3920 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3915(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3912(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3916(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3915 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3912 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3907(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3904(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3908(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3907 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3904 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3899(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3896(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3900(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3899 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3896 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3891(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3888(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3892(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3891 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3888 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3883(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3880(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3884(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3883 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3880 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3875(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3872(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3876(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3875 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3872 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3867(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3864(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3868(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3867 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3864 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3859(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3856(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3860(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3859 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3856 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3851(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3848(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3852(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3851 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3848 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3843(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3840(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3844(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3843 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3840 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3835(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3832(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3836(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3835 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3832 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3827(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3824(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3828(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3827 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3824 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3819(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3816(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3820(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3819 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3816 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3811(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3808(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3812(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3811 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3808 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3803(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3800(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3804(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3803 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3800 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3795(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3792(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3796(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3795 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3792 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3787(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3784(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3788(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3787 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3784 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3779(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3776(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3780(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3779 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3776 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3771(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3768(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3772(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3771 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3768 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3763(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3760(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3764(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3763 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3760 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3755(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3752(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3756(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3755 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3752 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3747(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3744(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3748(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3747 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3744 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3739(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3736(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3740(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3739 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3736 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3731(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3728(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3732(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3731 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3728 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3723(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3720(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3724(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3723 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3720 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3715(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3712(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3716(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3715 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3712 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3707(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3704(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3708(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3707 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3704 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3699(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3696(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3700(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3699 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3696 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3691(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3688(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3692(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3691 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3688 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3683(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3680(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3684(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3683 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3680 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3675(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3672(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3676(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3675 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3672 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3667(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3664(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3668(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3667 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3664 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3659(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3656(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3660(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3659 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3656 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3651(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3648(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3652(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3651 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3648 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3643(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3640(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3644(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3643 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3640 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3635(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3632(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3636(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3635 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3632 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3627(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3624(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3628(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3627 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3624 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3619(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3616(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3620(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3619 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3616 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3611(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3608(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3612(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3611 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3608 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3603(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3600(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3604(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3603 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3600 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3595(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3592(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3596(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3595 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3592 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3587(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3584(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3588(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3587 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3584 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3579(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3576(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3580(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3579 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3576 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3571(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_3568(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_3572(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_3571 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_3568 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__1_3539(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3540(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_3539 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_3531(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3528(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3532(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3531 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3528 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3523(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3520(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3524(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3523 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3520 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3515(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3512(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3516(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3515 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3512 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3507(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3504(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3508(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3507 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3504 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3499(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3496(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3500(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3499 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3496 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3491(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3488(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3492(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3491 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3488 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3483(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3480(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3484(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3483 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3480 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3475(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3472(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3476(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3475 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3472 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3467(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3464(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3468(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3467 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3464 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3459(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3456(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3460(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3459 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3456 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3451(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3448(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3452(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3451 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3448 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3443(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3440(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3444(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3443 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3440 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3435(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3432(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3436(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3435 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3432 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3427(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3424(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3428(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3427 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3424 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3419(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3416(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3420(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3419 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3416 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3411(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3408(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3412(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3411 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3408 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3403(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3400(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3404(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3403 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3400 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3395(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3392(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3396(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3395 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3392 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3387(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3384(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3388(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3387 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3384 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3379(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3376(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3380(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3379 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3376 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3371(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3368(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3372(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3371 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3368 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3363(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3360(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3364(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3363 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3360 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3355(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3352(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3356(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3355 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3352 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3347(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3344(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3348(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3347 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3344 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3339(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3336(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3340(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3339 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3336 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3331(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3328(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3332(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3331 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3328 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3323(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3320(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3324(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3323 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3320 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3315(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3312(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3316(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3315 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3312 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3307(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3304(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3308(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3307 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3304 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3299(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3296(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3300(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3299 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3296 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3291(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3288(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3292(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3291 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3288 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3283(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3280(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3284(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3283 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3280 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3275(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3272(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3276(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3275 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3272 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3267(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3264(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3268(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3267 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3264 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3259(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3256(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3260(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3259 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3256 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3251(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3248(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3252(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3251 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3248 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3243(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3240(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3244(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3243 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3240 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3235(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3232(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3236(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3235 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3232 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3227(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3224(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3228(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3227 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3224 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3219(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3216(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3220(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3219 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3216 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3211(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3208(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3212(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3211 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3208 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3203(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3200(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3204(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3203 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3200 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3195(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3192(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3196(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3195 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3192 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3187(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3184(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3188(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3187 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3184 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3179(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3176(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3180(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3179 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3176 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3171(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3168(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3172(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3171 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3168 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3163(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3160(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3164(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3163 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3160 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3155(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3152(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3156(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3155 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3152 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3147(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3144(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3148(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3147 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3144 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3139(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3136(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3140(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3139 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3136 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3131(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3128(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3132(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3131 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3128 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3123(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3120(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3124(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3123 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3120 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3115(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3112(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3116(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3115 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3112 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3107(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3104(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3108(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3107 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3104 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3099(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3096(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3100(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3099 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3096 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3091(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3088(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3092(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3091 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3088 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3083(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_3080(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_3084(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_3083 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_3080 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_3075(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_3072(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_3076(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_3075 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_3072 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__1_4093(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__1_4044 genblk1_4_a (.a(x[4]), .b(y[4]), .cin(), .sum(s[4]), 
      .carry(c1[4]));
   fulladder__1_4036 genblk1_5_a (.a(x[5]), .b(y[5]), .cin(z[5]), .sum(s1[5]), 
      .carry(c1[5]));
   fulladder__1_4028 genblk1_6_a (.a(x[6]), .b(y[6]), .cin(z[6]), .sum(s1[6]), 
      .carry(c1[6]));
   fulladder__1_4020 genblk1_7_a (.a(x[7]), .b(y[7]), .cin(z[7]), .sum(s1[7]), 
      .carry(c1[7]));
   fulladder__1_4012 genblk1_8_a (.a(x[8]), .b(y[8]), .cin(z[8]), .sum(s1[8]), 
      .carry(c1[8]));
   fulladder__1_4004 genblk1_9_a (.a(x[9]), .b(y[9]), .cin(z[9]), .sum(s1[9]), 
      .carry(c1[9]));
   fulladder__1_3996 genblk1_10_a (.a(x[10]), .b(y[10]), .cin(z[10]), .sum(
      s1[10]), .carry(c1[10]));
   fulladder__1_3988 genblk1_11_a (.a(x[11]), .b(y[11]), .cin(z[11]), .sum(
      s1[11]), .carry(c1[11]));
   fulladder__1_3980 genblk1_12_a (.a(x[12]), .b(y[12]), .cin(z[12]), .sum(
      s1[12]), .carry(c1[12]));
   fulladder__1_3972 genblk1_13_a (.a(x[13]), .b(y[13]), .cin(z[13]), .sum(
      s1[13]), .carry(c1[13]));
   fulladder__1_3964 genblk1_14_a (.a(x[14]), .b(y[14]), .cin(z[14]), .sum(
      s1[14]), .carry(c1[14]));
   fulladder__1_3956 genblk1_15_a (.a(x[15]), .b(y[15]), .cin(z[15]), .sum(
      s1[15]), .carry(c1[15]));
   fulladder__1_3948 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(z[16]), .sum(
      s1[16]), .carry(c1[16]));
   fulladder__1_3940 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(z[17]), .sum(
      s1[17]), .carry(c1[17]));
   fulladder__1_3932 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(
      s1[18]), .carry(c1[18]));
   fulladder__1_3924 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(
      s1[19]), .carry(c1[19]));
   fulladder__1_3916 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(
      s1[20]), .carry(c1[20]));
   fulladder__1_3908 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(
      s1[21]), .carry(c1[21]));
   fulladder__1_3900 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(
      s1[22]), .carry(c1[22]));
   fulladder__1_3892 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__1_3884 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__1_3876 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__1_3868 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__1_3860 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__1_3852 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__1_3844 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__1_3836 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__1_3828 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__1_3820 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__1_3812 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__1_3804 genblk1_34_a (.a(x[63]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__1_3796 genblk1_35_a (.a(x[63]), .b(y[63]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__1_3788 genblk1_36_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__1_3780 genblk1_37_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__1_3772 genblk1_38_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__1_3764 genblk1_39_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__1_3756 genblk1_40_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__1_3748 genblk1_41_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__1_3740 genblk1_42_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__1_3732 genblk1_43_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__1_3724 genblk1_44_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__1_3716 genblk1_45_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__1_3708 genblk1_46_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__1_3700 genblk1_47_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__1_3692 genblk1_48_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__1_3684 genblk1_49_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__1_3676 genblk1_50_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__1_3668 genblk1_51_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__1_3660 genblk1_52_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__1_3652 genblk1_53_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__1_3644 genblk1_54_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__1_3636 genblk1_55_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__1_3628 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__1_3620 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__1_3612 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__1_3604 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__1_3596 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__1_3588 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__1_3580 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__1_3572 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__1_3540 genblk2_4_b (.a(s1[5]), .b(c1[4]), .cin(), .sum(s[5]), 
      .carry(c2[5]));
   fulladder__1_3532 genblk2_5_b (.a(s1[6]), .b(c1[5]), .cin(c2[5]), .sum(s[6]), 
      .carry(c2[6]));
   fulladder__1_3524 genblk2_6_b (.a(s1[7]), .b(c1[6]), .cin(c2[6]), .sum(s[7]), 
      .carry(c2[7]));
   fulladder__1_3516 genblk2_7_b (.a(s1[8]), .b(c1[7]), .cin(c2[7]), .sum(s[8]), 
      .carry(c2[8]));
   fulladder__1_3508 genblk2_8_b (.a(s1[9]), .b(c1[8]), .cin(c2[8]), .sum(s[9]), 
      .carry(c2[9]));
   fulladder__1_3500 genblk2_9_b (.a(s1[10]), .b(c1[9]), .cin(c2[9]), .sum(s[10]), 
      .carry(c2[10]));
   fulladder__1_3492 genblk2_10_b (.a(s1[11]), .b(c1[10]), .cin(c2[10]), 
      .sum(s[11]), .carry(c2[11]));
   fulladder__1_3484 genblk2_11_b (.a(s1[12]), .b(c1[11]), .cin(c2[11]), 
      .sum(s[12]), .carry(c2[12]));
   fulladder__1_3476 genblk2_12_b (.a(s1[13]), .b(c1[12]), .cin(c2[12]), 
      .sum(s[13]), .carry(c2[13]));
   fulladder__1_3468 genblk2_13_b (.a(s1[14]), .b(c1[13]), .cin(c2[13]), 
      .sum(s[14]), .carry(c2[14]));
   fulladder__1_3460 genblk2_14_b (.a(s1[15]), .b(c1[14]), .cin(c2[14]), 
      .sum(s[15]), .carry(c2[15]));
   fulladder__1_3452 genblk2_15_b (.a(s1[16]), .b(c1[15]), .cin(c2[15]), 
      .sum(s[16]), .carry(c2[16]));
   fulladder__1_3444 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(c2[16]), 
      .sum(s[17]), .carry(c2[17]));
   fulladder__1_3436 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), 
      .sum(s[18]), .carry(c2[18]));
   fulladder__1_3428 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), 
      .sum(s[19]), .carry(c2[19]));
   fulladder__1_3420 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), 
      .sum(s[20]), .carry(c2[20]));
   fulladder__1_3412 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), 
      .sum(s[21]), .carry(c2[21]));
   fulladder__1_3404 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), 
      .sum(s[22]), .carry(c2[22]));
   fulladder__1_3396 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), 
      .sum(s[23]), .carry(c2[23]));
   fulladder__1_3388 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__1_3380 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__1_3372 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__1_3364 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__1_3356 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__1_3348 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__1_3340 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__1_3332 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__1_3324 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__1_3316 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__1_3308 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__1_3300 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__1_3292 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__1_3284 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__1_3276 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__1_3268 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__1_3260 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__1_3252 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__1_3244 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__1_3236 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__1_3228 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__1_3220 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__1_3212 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__1_3204 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__1_3196 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__1_3188 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__1_3180 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__1_3172 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__1_3164 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__1_3156 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__1_3148 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__1_3140 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__1_3132 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__1_3124 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__1_3116 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__1_3108 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__1_3100 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__1_3092 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__1_3084 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__1_3076 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__1_5044(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5045(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_5044 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_5036(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5033(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5037(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5036 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5033 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5028(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5025(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5029(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5028 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5025 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5020(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5017(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5021(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5020 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5017 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5012(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5009(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5013(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5012 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5009 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5004(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5001(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5005(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5004 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5001 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4996(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4993(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4997(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4996 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4993 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4988(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4985(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4989(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4988 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4985 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4980(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4977(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4981(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4980 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4977 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4972(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4969(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4973(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4972 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4969 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4964(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4961(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4965(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4964 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4961 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4956(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4953(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4957(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4956 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4953 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4948(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4945(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4949(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4948 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4945 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4940(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4937(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4941(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4940 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4937 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4932(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4929(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4933(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4932 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4929 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4924(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4921(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4925(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4924 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4921 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4916(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4913(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4917(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4916 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4913 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4908(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4905(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4909(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4908 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4905 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4900(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4897(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4901(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4900 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4897 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4892(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4889(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4893(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4892 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4889 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4884(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4881(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4885(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4884 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4881 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4876(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4873(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4877(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4876 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4873 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4868(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4865(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4869(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4868 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4865 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4860(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4857(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4861(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4860 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4857 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4852(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4849(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4853(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4852 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4849 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4844(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4841(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4845(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4844 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4841 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4836(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4833(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4837(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4836 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4833 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4828(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4825(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4829(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4828 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4825 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4820(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4817(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4821(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4820 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4817 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4812(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4809(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4813(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4812 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4809 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4804(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4801(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4805(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4804 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4801 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4796(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4793(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4797(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4796 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4793 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4788(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4789(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4788 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4785 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4780(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4781(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4780 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4777 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4772(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4773(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4772 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4769 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4764(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4765(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4764 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4761 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4756(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4757(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4756 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4753 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4748(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4745(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4749(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4748 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4745 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4740(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4737(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4741(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4740 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4737 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4732(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4729(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4733(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4732 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4729 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4724(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4721(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4725(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4724 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4721 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4716(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4713(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4717(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4716 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4713 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4708(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4705(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4709(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4708 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4705 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4700(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4697(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4701(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4700 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4697 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4692(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4689(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4693(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4692 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4689 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4684(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4681(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4685(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4684 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4681 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4676(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4673(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4677(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4676 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4673 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4668(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4665(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4669(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4668 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4665 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4660(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4657(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4661(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4660 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4657 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4652(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4649(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4653(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4652 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4649 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4644(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4641(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4645(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4644 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4641 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4636(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4633(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4637(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4636 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4633 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4628(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4625(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4629(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4628 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4625 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4620(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4617(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4621(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4620 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4617 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4612(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4609(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4613(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4612 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4609 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4604(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4601(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4605(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4604 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4601 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4596(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_4593(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_4597(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_4596 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_4593 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__1_4540(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4541(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_4540 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_4532(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4533(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4532 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4529 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4524(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4525(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4524 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4521 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4516(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4513(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4517(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4516 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4513 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4508(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4505(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4509(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4508 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4505 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4500(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4497(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4501(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4500 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4497 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4492(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4489(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4493(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4492 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4489 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4484(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4481(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4485(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4484 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4481 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4476(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4473(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4477(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4476 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4473 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4468(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4465(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4469(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4468 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4465 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4460(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4457(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4461(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4460 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4457 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4452(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4449(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4453(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4452 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4449 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4444(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4441(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4445(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4444 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4441 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4436(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4433(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4437(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4436 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4433 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4428(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4425(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4429(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4428 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4425 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4420(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4417(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4421(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4420 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4417 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4412(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4409(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4413(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4412 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4409 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4404(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4401(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4405(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4404 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4401 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4396(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4393(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4397(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4396 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4393 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4388(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4385(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4389(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4388 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4385 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4380(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4377(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4381(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4380 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4377 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4372(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4369(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4373(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4372 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4369 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4364(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4361(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4365(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4364 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4361 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4356(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4353(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4357(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4356 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4353 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4348(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4345(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4349(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4348 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4345 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4340(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4337(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4341(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4340 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4337 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4332(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4329(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4333(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4332 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4329 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4324(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4321(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4325(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4324 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4321 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4316(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4313(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4317(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4316 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4313 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4308(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4305(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4309(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4308 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4305 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4300(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4297(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4301(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4300 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4297 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4292(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4289(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4293(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4292 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4289 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4284(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4285(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4284 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4281 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4276(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4277(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4276 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4273 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4268(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4269(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4268 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4265 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4260(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4261(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4260 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4257 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4252(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4253(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4252 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4249 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4244(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4241(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4245(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4244 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4241 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4236(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4233(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4237(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4236 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4233 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4228(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4225(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4229(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4228 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4225 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4220(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4217(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4221(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4220 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4217 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4212(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4209(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4213(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4212 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4209 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4204(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4201(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4205(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4204 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4201 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4196(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4193(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4197(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4196 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4193 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4188(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4185(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4189(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4188 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4185 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4180(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4177(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4181(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4180 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4177 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4172(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4169(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4173(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4172 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4169 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4164(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4161(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4165(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4164 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4161 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4156(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4153(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4157(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4156 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4153 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4148(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4145(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4149(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4148 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4145 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4140(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4137(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4141(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4140 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4137 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4132(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4129(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4133(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4132 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4129 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4124(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4121(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4125(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4124 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4121 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4116(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4113(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4117(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4116 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4113 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4108(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_4105(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_4109(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_4108 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_4105 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_4100(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_4097(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_4101(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_4100 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_4097 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__1_5118(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__1_5045 genblk1_7_a (.a(x[7]), .b(y[7]), .cin(), .sum(s[7]), 
      .carry(c1[7]));
   fulladder__1_5037 genblk1_8_a (.a(x[8]), .b(y[8]), .cin(z[8]), .sum(s1[8]), 
      .carry(c1[8]));
   fulladder__1_5029 genblk1_9_a (.a(x[9]), .b(y[9]), .cin(z[9]), .sum(s1[9]), 
      .carry(c1[9]));
   fulladder__1_5021 genblk1_10_a (.a(x[10]), .b(y[10]), .cin(z[10]), .sum(
      s1[10]), .carry(c1[10]));
   fulladder__1_5013 genblk1_11_a (.a(x[11]), .b(y[11]), .cin(z[11]), .sum(
      s1[11]), .carry(c1[11]));
   fulladder__1_5005 genblk1_12_a (.a(x[12]), .b(y[12]), .cin(z[12]), .sum(
      s1[12]), .carry(c1[12]));
   fulladder__1_4997 genblk1_13_a (.a(x[13]), .b(y[13]), .cin(z[13]), .sum(
      s1[13]), .carry(c1[13]));
   fulladder__1_4989 genblk1_14_a (.a(x[14]), .b(y[14]), .cin(z[14]), .sum(
      s1[14]), .carry(c1[14]));
   fulladder__1_4981 genblk1_15_a (.a(x[15]), .b(y[15]), .cin(z[15]), .sum(
      s1[15]), .carry(c1[15]));
   fulladder__1_4973 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(z[16]), .sum(
      s1[16]), .carry(c1[16]));
   fulladder__1_4965 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(z[17]), .sum(
      s1[17]), .carry(c1[17]));
   fulladder__1_4957 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(
      s1[18]), .carry(c1[18]));
   fulladder__1_4949 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(
      s1[19]), .carry(c1[19]));
   fulladder__1_4941 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(
      s1[20]), .carry(c1[20]));
   fulladder__1_4933 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(
      s1[21]), .carry(c1[21]));
   fulladder__1_4925 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(
      s1[22]), .carry(c1[22]));
   fulladder__1_4917 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__1_4909 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__1_4901 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__1_4893 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__1_4885 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__1_4877 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__1_4869 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__1_4861 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__1_4853 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__1_4845 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__1_4837 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__1_4829 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__1_4821 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__1_4813 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__1_4805 genblk1_37_a (.a(x[63]), .b(y[37]), .cin(z[37]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__1_4797 genblk1_38_a (.a(x[63]), .b(y[63]), .cin(z[38]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__1_4789 genblk1_39_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__1_4781 genblk1_40_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__1_4773 genblk1_41_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__1_4765 genblk1_42_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__1_4757 genblk1_43_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__1_4749 genblk1_44_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__1_4741 genblk1_45_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__1_4733 genblk1_46_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__1_4725 genblk1_47_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__1_4717 genblk1_48_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__1_4709 genblk1_49_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__1_4701 genblk1_50_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__1_4693 genblk1_51_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__1_4685 genblk1_52_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__1_4677 genblk1_53_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__1_4669 genblk1_54_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__1_4661 genblk1_55_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__1_4653 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__1_4645 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__1_4637 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__1_4629 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__1_4621 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__1_4613 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__1_4605 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__1_4597 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__1_4541 genblk2_7_b (.a(s1[8]), .b(c1[7]), .cin(), .sum(s[8]), 
      .carry(c2[8]));
   fulladder__1_4533 genblk2_8_b (.a(s1[9]), .b(c1[8]), .cin(c2[8]), .sum(s[9]), 
      .carry(c2[9]));
   fulladder__1_4525 genblk2_9_b (.a(s1[10]), .b(c1[9]), .cin(c2[9]), .sum(s[10]), 
      .carry(c2[10]));
   fulladder__1_4517 genblk2_10_b (.a(s1[11]), .b(c1[10]), .cin(c2[10]), 
      .sum(s[11]), .carry(c2[11]));
   fulladder__1_4509 genblk2_11_b (.a(s1[12]), .b(c1[11]), .cin(c2[11]), 
      .sum(s[12]), .carry(c2[12]));
   fulladder__1_4501 genblk2_12_b (.a(s1[13]), .b(c1[12]), .cin(c2[12]), 
      .sum(s[13]), .carry(c2[13]));
   fulladder__1_4493 genblk2_13_b (.a(s1[14]), .b(c1[13]), .cin(c2[13]), 
      .sum(s[14]), .carry(c2[14]));
   fulladder__1_4485 genblk2_14_b (.a(s1[15]), .b(c1[14]), .cin(c2[14]), 
      .sum(s[15]), .carry(c2[15]));
   fulladder__1_4477 genblk2_15_b (.a(s1[16]), .b(c1[15]), .cin(c2[15]), 
      .sum(s[16]), .carry(c2[16]));
   fulladder__1_4469 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(c2[16]), 
      .sum(s[17]), .carry(c2[17]));
   fulladder__1_4461 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), 
      .sum(s[18]), .carry(c2[18]));
   fulladder__1_4453 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), 
      .sum(s[19]), .carry(c2[19]));
   fulladder__1_4445 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), 
      .sum(s[20]), .carry(c2[20]));
   fulladder__1_4437 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), 
      .sum(s[21]), .carry(c2[21]));
   fulladder__1_4429 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), 
      .sum(s[22]), .carry(c2[22]));
   fulladder__1_4421 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), 
      .sum(s[23]), .carry(c2[23]));
   fulladder__1_4413 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__1_4405 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__1_4397 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__1_4389 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__1_4381 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__1_4373 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__1_4365 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__1_4357 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__1_4349 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__1_4341 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__1_4333 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__1_4325 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__1_4317 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__1_4309 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__1_4301 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__1_4293 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__1_4285 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__1_4277 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__1_4269 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__1_4261 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__1_4253 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__1_4245 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__1_4237 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__1_4229 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__1_4221 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__1_4213 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__1_4205 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__1_4197 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__1_4189 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__1_4181 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__1_4173 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__1_4165 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__1_4157 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__1_4149 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__1_4141 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__1_4133 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__1_4125 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__1_4117 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__1_4109 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__1_4101 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__1_6029(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6030(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_6029 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_6021(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6022(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_6021 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_6013(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6014(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_6013 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_6005(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6002(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6006(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6005 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6002 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5997(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5994(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5998(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5997 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5994 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5989(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5986(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5990(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5989 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5986 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5981(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5978(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5982(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5981 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5978 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5973(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5970(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5974(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5973 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5970 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5965(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5962(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5966(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5965 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5962 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5957(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5954(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5958(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5957 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5954 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5949(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5946(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5950(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5949 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5946 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5941(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5938(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5942(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5941 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5938 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5933(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5930(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5934(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5933 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5930 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5925(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5922(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5926(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5925 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5922 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5917(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5914(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5918(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5917 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5914 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5909(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5906(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5910(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5909 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5906 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5901(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5898(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5902(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5901 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5898 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5893(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5890(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5894(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5893 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5890 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5885(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5882(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5886(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5885 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5882 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5877(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5874(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5878(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5877 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5874 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5869(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5866(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5870(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5869 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5866 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5861(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5858(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5862(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5861 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5858 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5853(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5850(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5854(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5853 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5850 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5845(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5842(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5846(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5845 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5842 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5837(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5834(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5838(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5837 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5834 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5829(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5826(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5830(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5829 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5826 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5821(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5818(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5822(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5821 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5818 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5813(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5810(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5814(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5813 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5810 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5805(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5802(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5806(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5805 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5802 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5797(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5794(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5798(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5797 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5794 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5789(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5786(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5790(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5789 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5786 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5781(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5778(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5782(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5781 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5778 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5773(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5770(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5774(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5773 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5770 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5765(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5762(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5766(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5765 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5762 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5757(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5754(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5758(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5757 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5754 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5749(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5746(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5750(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5749 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5746 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5741(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5738(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5742(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5741 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5738 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5733(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5730(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5734(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5733 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5730 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5725(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5722(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5726(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5725 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5722 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5717(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5714(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5718(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5717 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5714 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5709(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5706(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5710(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5709 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5706 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5701(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5698(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5702(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5701 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5698 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5693(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5690(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5694(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5693 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5690 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5685(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5682(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5686(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5685 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5682 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5677(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5674(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5678(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5677 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5674 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5669(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5666(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5670(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5669 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5666 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5661(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5658(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5662(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5661 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5658 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5653(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5650(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5654(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5653 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5650 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5645(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5642(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5646(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5645 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5642 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5637(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5634(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5638(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5637 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5634 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5629(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5626(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5630(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5629 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5626 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5621(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_5618(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_5622(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_5621 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_5618 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__1_5525(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5526(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_5525 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_5517(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5514(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5518(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5517 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5514 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5509(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5506(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5510(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5509 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5506 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5501(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5498(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5502(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5501 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5498 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5493(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5490(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5494(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5493 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5490 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5485(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5482(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5486(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5485 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5482 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5477(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5474(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5478(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5477 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5474 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5469(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5466(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5470(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5469 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5466 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5461(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5458(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5462(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5461 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5458 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5453(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5450(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5454(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5453 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5450 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5445(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5442(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5446(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5445 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5442 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5437(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5434(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5438(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5437 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5434 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5429(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5426(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5430(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5429 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5426 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5421(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5418(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5422(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5421 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5418 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5413(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5410(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5414(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5413 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5410 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5405(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5402(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5406(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5405 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5402 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5397(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5394(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5398(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5397 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5394 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5389(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5386(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5390(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5389 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5386 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5381(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5378(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5382(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5381 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5378 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5373(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5370(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5374(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5373 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5370 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5365(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5362(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5366(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5365 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5362 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5357(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5354(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5358(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5357 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5354 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5349(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5346(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5350(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5349 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5346 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5341(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5338(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5342(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5341 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5338 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5333(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5330(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5334(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5333 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5330 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5325(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5322(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5326(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5325 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5322 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5317(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5314(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5318(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5317 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5314 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5309(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5306(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5310(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5309 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5306 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5301(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5298(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5302(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5301 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5298 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5293(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5290(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5294(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5293 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5290 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5285(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5282(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5286(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5285 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5282 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5277(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5274(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5278(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5277 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5274 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5269(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5266(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5270(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5269 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5266 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5261(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5258(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5262(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5261 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5258 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5253(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5250(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5254(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5253 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5250 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5245(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5242(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5246(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5245 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5242 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5237(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5234(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5238(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5237 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5234 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5229(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5226(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5230(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5229 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5226 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5221(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5218(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5222(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5221 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5218 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5213(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5210(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5214(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5213 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5210 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5205(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5202(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5206(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5205 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5202 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5197(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5194(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5198(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5197 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5194 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5189(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5186(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5190(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5189 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5186 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5181(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5178(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5182(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5181 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5178 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5173(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5170(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5174(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5173 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5170 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5165(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5162(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5166(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5165 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5162 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5157(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5154(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5158(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5157 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5154 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5149(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5146(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5150(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5149 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5146 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5141(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5138(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5142(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5141 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5138 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5133(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_5130(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_5134(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_5133 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_5130 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_5125(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_5122(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_5126(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_5125 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_5122 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__1_6143(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__1_6030 genblk1_12_a (.a(x[12]), .b(y[12]), .cin(), .sum(s[12]), 
      .carry(c1[12]));
   fulladder__1_6022 genblk1_13_a (.a(x[13]), .b(y[13]), .cin(), .sum(s1[13]), 
      .carry(c1[13]));
   fulladder__1_6014 genblk1_14_a (.a(x[14]), .b(y[14]), .cin(), .sum(s1[14]), 
      .carry(c1[14]));
   fulladder__1_6006 genblk1_15_a (.a(x[15]), .b(y[15]), .cin(z[15]), .sum(
      s1[15]), .carry(c1[15]));
   fulladder__1_5998 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(z[16]), .sum(
      s1[16]), .carry(c1[16]));
   fulladder__1_5990 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(z[17]), .sum(
      s1[17]), .carry(c1[17]));
   fulladder__1_5982 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(
      s1[18]), .carry(c1[18]));
   fulladder__1_5974 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(
      s1[19]), .carry(c1[19]));
   fulladder__1_5966 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(
      s1[20]), .carry(c1[20]));
   fulladder__1_5958 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(
      s1[21]), .carry(c1[21]));
   fulladder__1_5950 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(
      s1[22]), .carry(c1[22]));
   fulladder__1_5942 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__1_5934 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__1_5926 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__1_5918 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__1_5910 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__1_5902 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__1_5894 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__1_5886 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__1_5878 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__1_5870 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__1_5862 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__1_5854 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__1_5846 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__1_5838 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__1_5830 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__1_5822 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__1_5814 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__1_5806 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__1_5798 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__1_5790 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__1_5782 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__1_5774 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__1_5766 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__1_5758 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__1_5750 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__1_5742 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__1_5734 genblk1_49_a (.a(x[49]), .b(y[49]), .cin(z[49]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__1_5726 genblk1_50_a (.a(x[50]), .b(y[50]), .cin(z[50]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__1_5718 genblk1_51_a (.a(x[51]), .b(y[51]), .cin(z[51]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__1_5710 genblk1_52_a (.a(x[52]), .b(y[52]), .cin(z[52]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__1_5702 genblk1_53_a (.a(x[53]), .b(y[53]), .cin(z[53]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__1_5694 genblk1_54_a (.a(x[54]), .b(y[54]), .cin(z[54]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__1_5686 genblk1_55_a (.a(x[55]), .b(y[55]), .cin(z[55]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__1_5678 genblk1_56_a (.a(x[56]), .b(y[56]), .cin(z[56]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__1_5670 genblk1_57_a (.a(x[57]), .b(y[57]), .cin(z[57]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__1_5662 genblk1_58_a (.a(x[58]), .b(y[58]), .cin(z[58]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__1_5654 genblk1_59_a (.a(x[59]), .b(y[59]), .cin(z[59]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__1_5646 genblk1_60_a (.a(x[60]), .b(y[60]), .cin(z[60]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__1_5638 genblk1_61_a (.a(x[61]), .b(y[61]), .cin(z[61]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__1_5630 genblk1_62_a (.a(x[62]), .b(y[62]), .cin(z[62]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__1_5622 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__1_5526 genblk2_12_b (.a(s1[13]), .b(c1[12]), .cin(), .sum(s[13]), 
      .carry(c2[13]));
   fulladder__1_5518 genblk2_13_b (.a(s1[14]), .b(c1[13]), .cin(c2[13]), 
      .sum(s[14]), .carry(c2[14]));
   fulladder__1_5510 genblk2_14_b (.a(s1[15]), .b(c1[14]), .cin(c2[14]), 
      .sum(s[15]), .carry(c2[15]));
   fulladder__1_5502 genblk2_15_b (.a(s1[16]), .b(c1[15]), .cin(c2[15]), 
      .sum(s[16]), .carry(c2[16]));
   fulladder__1_5494 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(c2[16]), 
      .sum(s[17]), .carry(c2[17]));
   fulladder__1_5486 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), 
      .sum(s[18]), .carry(c2[18]));
   fulladder__1_5478 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), 
      .sum(s[19]), .carry(c2[19]));
   fulladder__1_5470 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), 
      .sum(s[20]), .carry(c2[20]));
   fulladder__1_5462 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), 
      .sum(s[21]), .carry(c2[21]));
   fulladder__1_5454 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), 
      .sum(s[22]), .carry(c2[22]));
   fulladder__1_5446 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), 
      .sum(s[23]), .carry(c2[23]));
   fulladder__1_5438 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__1_5430 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__1_5422 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__1_5414 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__1_5406 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__1_5398 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__1_5390 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__1_5382 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__1_5374 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__1_5366 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__1_5358 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__1_5350 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__1_5342 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__1_5334 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__1_5326 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__1_5318 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__1_5310 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__1_5302 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__1_5294 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__1_5286 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__1_5278 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__1_5270 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__1_5262 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__1_5254 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__1_5246 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__1_5238 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__1_5230 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__1_5222 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__1_5214 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__1_5206 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__1_5198 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__1_5190 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__1_5182 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__1_5174 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__1_5166 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__1_5158 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__1_5150 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__1_5142 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__1_5134 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__1_5126 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__1_7070(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7071(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_7070 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_7062(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7059(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7063(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7062 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7059 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7054(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7051(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7055(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7054 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7051 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7046(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7043(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7047(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7046 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7043 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7038(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7035(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7039(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7038 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7035 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7030(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7027(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7031(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7030 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7027 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7022(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7019(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7023(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7022 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7019 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7014(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7011(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7015(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7014 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7011 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7006(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7003(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7007(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7006 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7003 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6998(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6995(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6999(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6998 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6995 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6990(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6987(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6991(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6990 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6987 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6982(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6979(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6983(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6982 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6979 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6974(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6971(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6975(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6974 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6971 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6966(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6963(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6967(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6966 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6963 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6958(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6955(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6959(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6958 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6955 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6950(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6947(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6951(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6950 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6947 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6942(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6939(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6943(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6942 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6939 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6934(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6931(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6935(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6934 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6931 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6926(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6923(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6927(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6926 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6923 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6918(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6915(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6919(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6918 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6915 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6910(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6907(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6911(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6910 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6907 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6902(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6899(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6903(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6902 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6899 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6894(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6891(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6895(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6894 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6891 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6886(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6883(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6887(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6886 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6883 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6878(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6875(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6879(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6878 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6875 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6870(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6867(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6871(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6870 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6867 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6862(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6859(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6863(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6862 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6859 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6854(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6851(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6855(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6854 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6851 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6846(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6843(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6847(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6846 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6843 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6838(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6835(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6839(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6838 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6835 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6830(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6827(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6831(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6830 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6827 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6822(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6819(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6823(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6822 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6819 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6814(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6811(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6815(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6814 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6811 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6806(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6803(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6807(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6806 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6803 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6798(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6795(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6799(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6798 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6795 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6790(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6787(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6791(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6790 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6787 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6782(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6779(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6783(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6782 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6779 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6771(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6775(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6774 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6771 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6763(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6767(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6766 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6763 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6755(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6759(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6758 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6755 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6750(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6747(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6751(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6750 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6747 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6742(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6739(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6743(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6742 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6739 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6734(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6731(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6735(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6734 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6731 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6726(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6723(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6727(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6726 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6723 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6718(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6715(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6719(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6718 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6715 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6710(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6707(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6711(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6710 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6707 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6702(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6699(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6703(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6702 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6699 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6694(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6691(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6695(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6694 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6691 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6686(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6683(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6687(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6686 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6683 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6678(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6675(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6679(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6678 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6675 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6670(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6667(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6671(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6670 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6667 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6662(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6659(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6663(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6662 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6659 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6654(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6651(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6655(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6654 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6651 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6646(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_6643(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_6647(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_6646 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_6643 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__1_6566(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6567(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_6566 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_6558(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6555(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6559(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6558 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6555 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6550(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6547(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6551(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6550 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6547 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6542(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6539(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6543(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6542 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6539 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6534(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6531(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6535(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6534 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6531 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6523(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6527(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6526 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6523 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6515(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6519(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6518 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6515 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6510(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6507(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6511(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6510 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6507 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6502(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6499(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6503(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6502 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6499 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6494(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6491(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6495(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6494 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6491 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6486(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6483(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6487(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6486 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6483 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6478(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6475(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6479(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6478 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6475 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6470(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6467(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6471(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6470 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6467 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6462(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6459(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6463(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6462 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6459 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6454(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6451(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6455(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6454 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6451 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6446(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6443(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6447(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6446 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6443 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6438(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6435(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6439(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6438 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6435 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6430(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6427(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6431(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6430 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6427 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6422(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6419(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6423(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6422 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6419 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6414(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6411(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6415(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6414 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6411 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6406(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6403(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6407(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6406 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6403 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6398(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6395(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6399(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6398 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6395 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6390(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6387(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6391(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6390 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6387 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6382(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6379(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6383(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6382 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6379 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6374(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6371(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6375(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6374 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6371 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6366(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6363(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6367(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6366 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6363 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6358(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6355(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6359(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6358 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6355 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6350(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6347(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6351(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6350 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6347 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6342(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6339(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6343(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6342 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6339 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6334(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6331(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6335(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6334 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6331 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6326(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6323(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6327(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6326 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6323 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6318(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6315(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6319(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6318 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6315 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6310(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6307(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6311(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6310 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6307 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6302(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6299(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6303(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6302 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6299 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6294(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6291(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6295(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6294 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6291 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6286(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6283(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6287(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6286 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6283 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6278(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6275(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6279(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6278 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6275 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6267(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6271(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6270 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6267 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6259(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6263(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6262 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6259 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6251(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6255(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6254 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6251 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6246(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6243(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6247(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6246 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6243 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6238(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6235(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6239(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6238 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6235 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6230(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6227(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6231(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6230 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6227 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6222(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6219(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6223(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6222 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6219 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6214(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6211(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6215(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6214 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6211 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6206(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6203(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6207(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6206 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6203 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6198(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6195(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6199(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6198 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6195 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6190(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6187(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6191(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6190 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6187 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6182(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6179(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6183(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6182 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6179 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6174(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6171(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6175(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6174 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6171 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6166(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6163(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6167(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6166 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6163 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6158(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_6155(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_6159(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_6158 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_6155 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_6150(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_6147(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_6151(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_6150 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_6147 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__1_7168(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__1_7071 genblk1_10_a (.a(x[10]), .b(y[10]), .cin(), .sum(s[10]), 
      .carry(c1[10]));
   fulladder__1_7063 genblk1_11_a (.a(x[11]), .b(y[11]), .cin(z[11]), .sum(
      s1[11]), .carry(c1[11]));
   fulladder__1_7055 genblk1_12_a (.a(x[12]), .b(y[12]), .cin(z[12]), .sum(
      s1[12]), .carry(c1[12]));
   fulladder__1_7047 genblk1_13_a (.a(x[13]), .b(y[13]), .cin(z[13]), .sum(
      s1[13]), .carry(c1[13]));
   fulladder__1_7039 genblk1_14_a (.a(x[14]), .b(y[14]), .cin(z[14]), .sum(
      s1[14]), .carry(c1[14]));
   fulladder__1_7031 genblk1_15_a (.a(x[15]), .b(y[15]), .cin(z[15]), .sum(
      s1[15]), .carry(c1[15]));
   fulladder__1_7023 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(z[16]), .sum(
      s1[16]), .carry(c1[16]));
   fulladder__1_7015 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(z[17]), .sum(
      s1[17]), .carry(c1[17]));
   fulladder__1_7007 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(
      s1[18]), .carry(c1[18]));
   fulladder__1_6999 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(
      s1[19]), .carry(c1[19]));
   fulladder__1_6991 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(
      s1[20]), .carry(c1[20]));
   fulladder__1_6983 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(
      s1[21]), .carry(c1[21]));
   fulladder__1_6975 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(
      s1[22]), .carry(c1[22]));
   fulladder__1_6967 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__1_6959 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__1_6951 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__1_6943 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__1_6935 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__1_6927 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__1_6919 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__1_6911 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__1_6903 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__1_6895 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__1_6887 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__1_6879 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__1_6871 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__1_6863 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__1_6855 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__1_6847 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__1_6839 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__1_6831 genblk1_40_a (.a(x[63]), .b(y[40]), .cin(z[40]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__1_6823 genblk1_41_a (.a(x[63]), .b(y[63]), .cin(z[41]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__1_6815 genblk1_42_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__1_6807 genblk1_43_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__1_6799 genblk1_44_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__1_6791 genblk1_45_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__1_6783 genblk1_46_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__1_6775 genblk1_47_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__1_6767 genblk1_48_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__1_6759 genblk1_49_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__1_6751 genblk1_50_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__1_6743 genblk1_51_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__1_6735 genblk1_52_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__1_6727 genblk1_53_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__1_6719 genblk1_54_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__1_6711 genblk1_55_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__1_6703 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__1_6695 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__1_6687 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__1_6679 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__1_6671 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__1_6663 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__1_6655 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__1_6647 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__1_6567 genblk2_10_b (.a(s1[11]), .b(c1[10]), .cin(), .sum(s[11]), 
      .carry(c2[11]));
   fulladder__1_6559 genblk2_11_b (.a(s1[12]), .b(c1[11]), .cin(c2[11]), 
      .sum(s[12]), .carry(c2[12]));
   fulladder__1_6551 genblk2_12_b (.a(s1[13]), .b(c1[12]), .cin(c2[12]), 
      .sum(s[13]), .carry(c2[13]));
   fulladder__1_6543 genblk2_13_b (.a(s1[14]), .b(c1[13]), .cin(c2[13]), 
      .sum(s[14]), .carry(c2[14]));
   fulladder__1_6535 genblk2_14_b (.a(s1[15]), .b(c1[14]), .cin(c2[14]), 
      .sum(s[15]), .carry(c2[15]));
   fulladder__1_6527 genblk2_15_b (.a(s1[16]), .b(c1[15]), .cin(c2[15]), 
      .sum(s[16]), .carry(c2[16]));
   fulladder__1_6519 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(c2[16]), 
      .sum(s[17]), .carry(c2[17]));
   fulladder__1_6511 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), 
      .sum(s[18]), .carry(c2[18]));
   fulladder__1_6503 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), 
      .sum(s[19]), .carry(c2[19]));
   fulladder__1_6495 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), 
      .sum(s[20]), .carry(c2[20]));
   fulladder__1_6487 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), 
      .sum(s[21]), .carry(c2[21]));
   fulladder__1_6479 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), 
      .sum(s[22]), .carry(c2[22]));
   fulladder__1_6471 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), 
      .sum(s[23]), .carry(c2[23]));
   fulladder__1_6463 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__1_6455 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__1_6447 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__1_6439 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__1_6431 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__1_6423 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__1_6415 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__1_6407 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__1_6399 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__1_6391 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__1_6383 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__1_6375 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__1_6367 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__1_6359 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__1_6351 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__1_6343 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__1_6335 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__1_6327 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__1_6319 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__1_6311 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__1_6303 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__1_6295 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__1_6287 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__1_6279 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__1_6271 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__1_6263 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__1_6255 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__1_6247 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__1_6239 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__1_6231 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__1_6223 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__1_6215 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__1_6207 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__1_6199 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__1_6191 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__1_6183 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__1_6175 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__1_6167 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__1_6159 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__1_6151 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__1_8071(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8072(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_8071 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_8063(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_8060(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8064(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_8063 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_8060 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_8055(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_8052(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8056(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_8055 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_8052 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_8047(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_8044(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8048(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_8047 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_8044 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_8039(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_8036(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8040(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_8039 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_8036 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_8031(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_8028(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8032(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_8031 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_8028 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_8023(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_8020(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8024(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_8023 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_8020 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_8015(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_8012(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8016(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_8015 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_8012 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_8007(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_8004(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8008(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_8007 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_8004 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7999(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7996(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_8000(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7999 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7996 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7991(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7988(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7992(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7991 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7988 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7983(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7980(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7984(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7983 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7980 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7975(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7972(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7976(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7975 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7972 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7967(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7964(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7968(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7967 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7964 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7959(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7956(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7960(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7959 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7956 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7951(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7948(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7952(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7951 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7948 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7943(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7940(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7944(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7943 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7940 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7935(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7932(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7936(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7935 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7932 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7927(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7924(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7928(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7927 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7924 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7919(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7916(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7920(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7919 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7916 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7911(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7908(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7912(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7911 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7908 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7903(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7900(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7904(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7903 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7900 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7895(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7892(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7896(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7895 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7892 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7887(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7884(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7888(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7887 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7884 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7879(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7876(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7880(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7879 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7876 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7871(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7868(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7872(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7871 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7868 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7863(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7860(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7864(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7863 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7860 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7855(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7852(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7856(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7855 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7852 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7847(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7844(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7848(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7847 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7844 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7839(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7836(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7840(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7839 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7836 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7831(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7828(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7832(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7831 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7828 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7823(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7820(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7824(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7823 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7820 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7815(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7812(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7816(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7815 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7812 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7807(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7804(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7808(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7807 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7804 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7799(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7796(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7800(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7799 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7796 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7791(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7788(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7792(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7791 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7788 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7783(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7780(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7784(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7783 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7780 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7775(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7772(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7776(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7775 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7772 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7767(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7764(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7768(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7767 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7764 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7759(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7756(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7760(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7759 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7756 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7751(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7748(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7752(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7751 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7748 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7743(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7740(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7744(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7743 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7740 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7735(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7732(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7736(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7735 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7732 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7727(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7724(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7728(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7727 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7724 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7719(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7716(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7720(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7719 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7716 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7711(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7708(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7712(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7711 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7708 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7703(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7700(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7704(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7703 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7700 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7695(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7692(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7696(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7695 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7692 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7687(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7684(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7688(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7687 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7684 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7679(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7676(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7680(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7679 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7676 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7671(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_7668(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_7672(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_7671 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_7668 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__1_7567(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7568(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_7567 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_7559(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7556(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7560(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7559 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7556 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7551(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7548(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7552(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7551 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7548 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7543(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7540(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7544(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7543 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7540 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7535(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7532(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7536(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7535 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7532 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7527(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7524(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7528(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7527 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7524 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7519(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7516(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7520(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7519 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7516 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7511(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7508(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7512(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7511 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7508 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7503(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7500(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7504(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7503 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7500 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7495(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7492(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7496(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7495 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7492 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7487(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7484(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7488(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7487 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7484 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7479(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7476(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7480(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7479 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7476 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7471(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7468(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7472(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7471 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7468 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7463(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7460(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7464(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7463 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7460 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7455(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7452(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7456(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7455 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7452 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7447(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7444(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7448(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7447 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7444 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7439(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7436(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7440(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7439 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7436 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7431(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7428(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7432(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7431 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7428 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7423(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7420(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7424(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7423 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7420 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7415(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7412(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7416(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7415 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7412 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7407(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7404(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7408(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7407 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7404 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7399(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7396(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7400(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7399 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7396 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7391(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7388(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7392(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7391 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7388 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7383(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7380(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7384(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7383 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7380 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7375(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7372(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7376(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7375 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7372 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7367(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7364(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7368(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7367 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7364 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7359(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7356(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7360(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7359 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7356 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7351(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7348(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7352(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7351 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7348 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7343(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7340(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7344(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7343 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7340 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7335(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7332(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7336(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7335 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7332 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7327(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7324(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7328(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7327 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7324 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7319(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7316(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7320(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7319 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7316 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7311(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7308(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7312(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7311 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7308 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7303(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7300(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7304(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7303 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7300 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7295(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7292(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7296(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7295 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7292 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7287(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7284(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7288(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7287 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7284 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7279(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7276(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7280(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7279 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7276 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7271(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7268(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7272(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7271 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7268 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7263(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7260(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7264(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7263 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7260 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7255(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7252(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7256(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7255 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7252 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7247(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7244(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7248(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7247 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7244 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7239(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7236(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7240(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7239 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7236 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7231(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7228(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7232(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7231 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7228 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7223(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7220(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7224(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7223 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7220 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7215(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7212(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7216(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7215 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7212 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7207(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7204(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7208(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7207 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7204 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7199(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7196(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7200(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7199 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7196 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7191(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7188(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7192(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7191 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7188 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7183(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_7180(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_7184(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_7183 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_7180 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_7175(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_7172(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_7176(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_7175 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_7172 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__1_8193(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__1_8072 genblk1_13_a (.a(x[13]), .b(y[13]), .cin(), .sum(s[13]), 
      .carry(c1[13]));
   fulladder__1_8064 genblk1_14_a (.a(x[14]), .b(y[14]), .cin(z[14]), .sum(
      s1[14]), .carry(c1[14]));
   fulladder__1_8056 genblk1_15_a (.a(x[15]), .b(y[15]), .cin(z[15]), .sum(
      s1[15]), .carry(c1[15]));
   fulladder__1_8048 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(z[16]), .sum(
      s1[16]), .carry(c1[16]));
   fulladder__1_8040 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(z[17]), .sum(
      s1[17]), .carry(c1[17]));
   fulladder__1_8032 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(
      s1[18]), .carry(c1[18]));
   fulladder__1_8024 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(
      s1[19]), .carry(c1[19]));
   fulladder__1_8016 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(
      s1[20]), .carry(c1[20]));
   fulladder__1_8008 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(
      s1[21]), .carry(c1[21]));
   fulladder__1_8000 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(
      s1[22]), .carry(c1[22]));
   fulladder__1_7992 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__1_7984 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__1_7976 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__1_7968 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__1_7960 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__1_7952 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__1_7944 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__1_7936 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__1_7928 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__1_7920 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__1_7912 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__1_7904 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__1_7896 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__1_7888 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__1_7880 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__1_7872 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__1_7864 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__1_7856 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__1_7848 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__1_7840 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__1_7832 genblk1_43_a (.a(x[63]), .b(y[43]), .cin(z[43]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__1_7824 genblk1_44_a (.a(x[63]), .b(y[63]), .cin(z[44]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__1_7816 genblk1_45_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__1_7808 genblk1_46_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__1_7800 genblk1_47_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__1_7792 genblk1_48_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__1_7784 genblk1_49_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__1_7776 genblk1_50_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__1_7768 genblk1_51_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__1_7760 genblk1_52_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__1_7752 genblk1_53_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__1_7744 genblk1_54_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__1_7736 genblk1_55_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__1_7728 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__1_7720 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__1_7712 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__1_7704 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__1_7696 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__1_7688 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__1_7680 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__1_7672 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__1_7568 genblk2_13_b (.a(s1[14]), .b(c1[13]), .cin(), .sum(s[14]), 
      .carry(c2[14]));
   fulladder__1_7560 genblk2_14_b (.a(s1[15]), .b(c1[14]), .cin(c2[14]), 
      .sum(s[15]), .carry(c2[15]));
   fulladder__1_7552 genblk2_15_b (.a(s1[16]), .b(c1[15]), .cin(c2[15]), 
      .sum(s[16]), .carry(c2[16]));
   fulladder__1_7544 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(c2[16]), 
      .sum(s[17]), .carry(c2[17]));
   fulladder__1_7536 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), 
      .sum(s[18]), .carry(c2[18]));
   fulladder__1_7528 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), 
      .sum(s[19]), .carry(c2[19]));
   fulladder__1_7520 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), 
      .sum(s[20]), .carry(c2[20]));
   fulladder__1_7512 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), 
      .sum(s[21]), .carry(c2[21]));
   fulladder__1_7504 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), 
      .sum(s[22]), .carry(c2[22]));
   fulladder__1_7496 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), 
      .sum(s[23]), .carry(c2[23]));
   fulladder__1_7488 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__1_7480 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__1_7472 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__1_7464 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__1_7456 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__1_7448 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__1_7440 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__1_7432 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__1_7424 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__1_7416 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__1_7408 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__1_7400 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__1_7392 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__1_7384 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__1_7376 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__1_7368 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__1_7360 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__1_7352 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__1_7344 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__1_7336 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__1_7328 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__1_7320 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__1_7312 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__1_7304 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__1_7296 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__1_7288 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__1_7280 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__1_7272 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__1_7264 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__1_7256 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__1_7248 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__1_7240 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__1_7232 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__1_7224 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__1_7216 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__1_7208 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__1_7200 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__1_7192 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__1_7184 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__1_7176 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__1_153(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_154(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_153 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_161(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_158(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_162(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_161 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_158 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_169(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_166(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_170(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_169 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_166 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_177(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_174(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_178(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_177 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_174 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_185(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_182(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_186(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_185 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_182 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_193(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_190(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_194(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_193 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_190 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_201(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_198(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_202(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_201 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_198 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_209(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_206(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_210(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_209 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_206 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_217(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_214(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_217 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_214 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_225(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_222(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_226(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_225 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_222 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_233(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_230(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_234(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_233 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_230 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_241(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_238(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_241 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_238 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_246(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_249 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_246 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_258(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_257 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_254 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_265 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_262 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_273 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_270 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_278(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_281 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_278 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_289(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_286(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_289 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_286 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_297(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_294(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_298(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_297 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_294 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_305(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_302(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_306(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_305 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_302 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_313(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_310(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_313 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_310 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_321(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_318(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_322(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_321 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_318 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_329(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_326(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_330(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_329 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_326 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_337(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_334(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_337 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_334 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_345(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_342(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_346(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_345 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_342 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_353(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_350(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_354(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_353 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_350 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_361(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_358(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_362(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_361 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_358 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_369(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_366(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_370(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_369 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_366 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_377(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_374(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_378(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_377 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_374 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_385(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_382(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_386(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_385 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_382 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_393(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_390(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_394(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_393 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_390 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_401(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_398(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_402(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_401 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_398 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_409(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_406(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_410(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_409 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_406 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_417(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_414(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_418(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_417 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_414 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_425(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_422(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_426(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_425 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_422 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_433(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_430(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_434(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_433 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_430 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_441(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_438(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_442(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_441 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_438 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_449(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_446(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_450(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_449 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_446 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_457(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_454(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_458(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_457 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_454 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_465(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_462(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_466(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_465 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_462 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_473(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_470(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_474(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_473 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_470 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_481(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_478(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_482(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_481 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_478 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_489(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_486(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_490(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_489 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_486 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_497(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_494(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_498(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_497 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_494 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_505(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_502(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_506(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_505 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_502 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_513(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_510(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_514(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_513 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_510 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_521 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_518 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__1_526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__1_530(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_529 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__1_526 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__1_657(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_658(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__1_657 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__1_665(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_662(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_666(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_665 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_662 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_673(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_670(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_674(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_673 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_670 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_681(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_678(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_682(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_681 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_678 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_689(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_686(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_690(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_689 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_686 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_697(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_694(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_698(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_697 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_694 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_705(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_702(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_706(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_705 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_702 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_713(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_710(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_714(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_713 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_710 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_721(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_718(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_722(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_721 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_718 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_729(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_726(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_730(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_729 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_726 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_737(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_734(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_737 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_734 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_745(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_742(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_745 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_742 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_750(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_753 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_750 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_761 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_758 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_769 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_766 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_778(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_777 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_774 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_782(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_785 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_782 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_793(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_790(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_793 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_790 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_801(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_798(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_802(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_801 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_798 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_809(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_806(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_809 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_806 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_817(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_814(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_817 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_814 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_825(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_822(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_826(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_825 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_822 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_833(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_830(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_833 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_830 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_841(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_838(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_842(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_841 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_838 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_849(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_846(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_850(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_849 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_846 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_857(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_854(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_858(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_857 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_854 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_865(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_862(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_866(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_865 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_862 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_873(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_870(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_874(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_873 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_870 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_881(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_878(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_882(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_881 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_878 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_889(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_886(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_890(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_889 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_886 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_897(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_894(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_898(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_897 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_894 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_905(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_902(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_906(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_905 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_902 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_913(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_910(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_914(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_913 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_910 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_921(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_918(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_922(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_921 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_918 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_929(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_926(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_930(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_929 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_926 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_937(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_934(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_938(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_937 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_934 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_945(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_942(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_946(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_945 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_942 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_953(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_950(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_954(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_953 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_950 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_961(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_958(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_962(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_961 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_958 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_969(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_966(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_970(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_969 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_966 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_977(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_974(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_978(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_977 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_974 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_985(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_982(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_986(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_985 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_982 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_993(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_990(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_994(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_993 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_990 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1001(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_998(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1002(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1001 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_998 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1009(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1006(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1010(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1009 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1006 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_1017(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__1_1014(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__1_1018(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__1_1017 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__1_1014 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__1_2(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__0_110(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__0_111(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__1_2 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__0_110 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__0_112(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__1_154 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(), .sum(s[16]), 
      .carry(c1[16]));
   fulladder__1_162 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(z[17]), .sum(s1[17]), 
      .carry(c1[17]));
   fulladder__1_170 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(s1[18]), 
      .carry(c1[18]));
   fulladder__1_178 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(s1[19]), 
      .carry(c1[19]));
   fulladder__1_186 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(s1[20]), 
      .carry(c1[20]));
   fulladder__1_194 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(s1[21]), 
      .carry(c1[21]));
   fulladder__1_202 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(s1[22]), 
      .carry(c1[22]));
   fulladder__1_210 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(s1[23]), 
      .carry(c1[23]));
   fulladder__1_218 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(s1[24]), 
      .carry(c1[24]));
   fulladder__1_226 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(s1[25]), 
      .carry(c1[25]));
   fulladder__1_234 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(s1[26]), 
      .carry(c1[26]));
   fulladder__1_242 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(s1[27]), 
      .carry(c1[27]));
   fulladder__1_250 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(s1[28]), 
      .carry(c1[28]));
   fulladder__1_258 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(s1[29]), 
      .carry(c1[29]));
   fulladder__1_266 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(s1[30]), 
      .carry(c1[30]));
   fulladder__1_274 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(s1[31]), 
      .carry(c1[31]));
   fulladder__1_282 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(s1[32]), 
      .carry(c1[32]));
   fulladder__1_290 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(s1[33]), 
      .carry(c1[33]));
   fulladder__1_298 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(s1[34]), 
      .carry(c1[34]));
   fulladder__1_306 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(s1[35]), 
      .carry(c1[35]));
   fulladder__1_314 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(s1[36]), 
      .carry(c1[36]));
   fulladder__1_322 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(s1[37]), 
      .carry(c1[37]));
   fulladder__1_330 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(s1[38]), 
      .carry(c1[38]));
   fulladder__1_338 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(s1[39]), 
      .carry(c1[39]));
   fulladder__1_346 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(s1[40]), 
      .carry(c1[40]));
   fulladder__1_354 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(s1[41]), 
      .carry(c1[41]));
   fulladder__1_362 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(s1[42]), 
      .carry(c1[42]));
   fulladder__1_370 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(s1[43]), 
      .carry(c1[43]));
   fulladder__1_378 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(s1[44]), 
      .carry(c1[44]));
   fulladder__1_386 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(s1[45]), 
      .carry(c1[45]));
   fulladder__1_394 genblk1_46_a (.a(x[63]), .b(y[46]), .cin(z[46]), .sum(s1[46]), 
      .carry(c1[46]));
   fulladder__1_402 genblk1_47_a (.a(x[63]), .b(y[63]), .cin(z[47]), .sum(s1[47]), 
      .carry(c1[47]));
   fulladder__1_410 genblk1_48_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[48]), 
      .carry(c1[48]));
   fulladder__1_418 genblk1_49_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[49]), 
      .carry(c1[49]));
   fulladder__1_426 genblk1_50_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[50]), 
      .carry(c1[50]));
   fulladder__1_434 genblk1_51_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[51]), 
      .carry(c1[51]));
   fulladder__1_442 genblk1_52_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[52]), 
      .carry(c1[52]));
   fulladder__1_450 genblk1_53_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[53]), 
      .carry(c1[53]));
   fulladder__1_458 genblk1_54_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[54]), 
      .carry(c1[54]));
   fulladder__1_466 genblk1_55_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[55]), 
      .carry(c1[55]));
   fulladder__1_474 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[56]), 
      .carry(c1[56]));
   fulladder__1_482 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[57]), 
      .carry(c1[57]));
   fulladder__1_490 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[58]), 
      .carry(c1[58]));
   fulladder__1_498 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[59]), 
      .carry(c1[59]));
   fulladder__1_506 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[60]), 
      .carry(c1[60]));
   fulladder__1_514 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[61]), 
      .carry(c1[61]));
   fulladder__1_522 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[62]), 
      .carry(c1[62]));
   fulladder__1_530 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[63]), 
      .carry());
   fulladder__1_658 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(), .sum(s[17]), 
      .carry(c2[17]));
   fulladder__1_666 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), .sum(
      s[18]), .carry(c2[18]));
   fulladder__1_674 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), .sum(
      s[19]), .carry(c2[19]));
   fulladder__1_682 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), .sum(
      s[20]), .carry(c2[20]));
   fulladder__1_690 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), .sum(
      s[21]), .carry(c2[21]));
   fulladder__1_698 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), .sum(
      s[22]), .carry(c2[22]));
   fulladder__1_706 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), .sum(
      s[23]), .carry(c2[23]));
   fulladder__1_714 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), .sum(
      s[24]), .carry(c2[24]));
   fulladder__1_722 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), .sum(
      s[25]), .carry(c2[25]));
   fulladder__1_730 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), .sum(
      s[26]), .carry(c2[26]));
   fulladder__1_738 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), .sum(
      s[27]), .carry(c2[27]));
   fulladder__1_746 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), .sum(
      s[28]), .carry(c2[28]));
   fulladder__1_754 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), .sum(
      s[29]), .carry(c2[29]));
   fulladder__1_762 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), .sum(
      s[30]), .carry(c2[30]));
   fulladder__1_770 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), .sum(
      s[31]), .carry(c2[31]));
   fulladder__1_778 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), .sum(
      s[32]), .carry(c2[32]));
   fulladder__1_786 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), .sum(
      s[33]), .carry(c2[33]));
   fulladder__1_794 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), .sum(
      s[34]), .carry(c2[34]));
   fulladder__1_802 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), .sum(
      s[35]), .carry(c2[35]));
   fulladder__1_810 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), .sum(
      s[36]), .carry(c2[36]));
   fulladder__1_818 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), .sum(
      s[37]), .carry(c2[37]));
   fulladder__1_826 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), .sum(
      s[38]), .carry(c2[38]));
   fulladder__1_834 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), .sum(
      s[39]), .carry(c2[39]));
   fulladder__1_842 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), .sum(
      s[40]), .carry(c2[40]));
   fulladder__1_850 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), .sum(
      s[41]), .carry(c2[41]));
   fulladder__1_858 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), .sum(
      s[42]), .carry(c2[42]));
   fulladder__1_866 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), .sum(
      s[43]), .carry(c2[43]));
   fulladder__1_874 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), .sum(
      s[44]), .carry(c2[44]));
   fulladder__1_882 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), .sum(
      s[45]), .carry(c2[45]));
   fulladder__1_890 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), .sum(
      s[46]), .carry(c2[46]));
   fulladder__1_898 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), .sum(
      s[47]), .carry(c2[47]));
   fulladder__1_906 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), .sum(
      s[48]), .carry(c2[48]));
   fulladder__1_914 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), .sum(
      s[49]), .carry(c2[49]));
   fulladder__1_922 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), .sum(
      s[50]), .carry(c2[50]));
   fulladder__1_930 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), .sum(
      s[51]), .carry(c2[51]));
   fulladder__1_938 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), .sum(
      s[52]), .carry(c2[52]));
   fulladder__1_946 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), .sum(
      s[53]), .carry(c2[53]));
   fulladder__1_954 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), .sum(
      s[54]), .carry(c2[54]));
   fulladder__1_962 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), .sum(
      s[55]), .carry(c2[55]));
   fulladder__1_970 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), .sum(
      s[56]), .carry(c2[56]));
   fulladder__1_978 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), .sum(
      s[57]), .carry(c2[57]));
   fulladder__1_986 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), .sum(
      s[58]), .carry(c2[58]));
   fulladder__1_994 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), .sum(
      s[59]), .carry(c2[59]));
   fulladder__1_1002 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__1_1010 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__1_1018 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__0_111 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), .sum(
      s[63]), .carry());
endmodule

module halfadder__2_49(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_50(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__2_49 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__2_57(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_58(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__2_57 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__2_65(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_66(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__2_65 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__2_73(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_70(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_74(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_73 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_70 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_81(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_78(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_82(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_81 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_78 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_89(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_86(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_90(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_89 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_86 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_97(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_94(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_98(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_97 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_94 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_105(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_102(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_106(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_105 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_102 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_113(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_110(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_114(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_113 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_110 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_121(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_118(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_122(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_121 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_118 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_129(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_126(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_130(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_129 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_126 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_137(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_134(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_138(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_137 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_134 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_145(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_142(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_146(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_145 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_142 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_153(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_150(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_154(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_153 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_150 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_161(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_158(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_162(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_161 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_158 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_169(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_166(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_170(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_169 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_166 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_177(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_174(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_178(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_177 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_174 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_185(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_182(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_186(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_185 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_182 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_193(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_190(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_194(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_193 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_190 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_201(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_198(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_202(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_201 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_198 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_209(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_206(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_210(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_209 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_206 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_217(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_214(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_217 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_214 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_225(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_222(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_226(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_225 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_222 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_233(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_230(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_234(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_233 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_230 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_241(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_238(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_241 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_238 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_246(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_249 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_246 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_258(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_257 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_254 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_265 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_262 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_273 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_270 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_278(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_281 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_278 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_289(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_286(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_289 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_286 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_297(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_294(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_298(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_297 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_294 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_305(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_302(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_306(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_305 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_302 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_313(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_310(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_313 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_310 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_321(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_318(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_322(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_321 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_318 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_329(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_326(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_330(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_329 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_326 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_337(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_334(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_337 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_334 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_345(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_342(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_346(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_345 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_342 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_353(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_350(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_354(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_353 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_350 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_361(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_358(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_362(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_361 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_358 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_369(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_366(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_370(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_369 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_366 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_377(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_374(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_378(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_377 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_374 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_385(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_382(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_386(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_385 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_382 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_393(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_390(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_394(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_393 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_390 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_401(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_398(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_402(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_401 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_398 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_409(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_406(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_410(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_409 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_406 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_417(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_414(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_418(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_417 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_414 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_425(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_422(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_426(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_425 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_422 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_433(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_430(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_434(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_433 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_430 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_441(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_438(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_442(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_441 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_438 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_449(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_446(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_450(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_449 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_446 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_457(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_454(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_458(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_457 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_454 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_465(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_462(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_466(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_465 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_462 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_473(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_470(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_474(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_473 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_470 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_481(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_478(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_482(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_481 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_478 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_489(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_486(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_490(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_489 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_486 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_497(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_494(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_498(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_497 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_494 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_505(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_502(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_506(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_505 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_502 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_513(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_510(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_514(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_513 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_510 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_521 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_518 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__2_526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__2_530(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__2_529 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__2_526 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__2_553(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_554(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__2_553 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__2_561(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_558(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_562(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_561 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_558 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_569(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_566(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_570(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_569 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_566 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_577(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_574(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_578(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_577 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_574 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_585(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_582(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_586(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_585 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_582 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_593(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_590(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_594(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_593 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_590 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_601(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_598(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_602(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_601 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_598 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_609(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_606(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_610(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_609 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_606 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_617(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_614(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_618(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_617 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_614 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_625(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_622(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_626(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_625 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_622 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_633(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_630(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_634(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_633 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_630 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_641(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_638(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_642(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_641 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_638 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_649(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_646(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_650(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_649 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_646 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_657(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_654(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_658(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_657 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_654 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_665(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_662(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_666(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_665 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_662 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_673(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_670(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_674(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_673 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_670 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_681(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_678(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_682(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_681 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_678 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_689(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_686(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_690(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_689 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_686 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_697(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_694(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_698(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_697 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_694 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_705(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_702(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_706(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_705 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_702 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_713(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_710(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_714(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_713 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_710 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_721(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_718(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_722(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_721 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_718 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_729(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_726(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_730(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_729 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_726 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_737(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_734(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_737 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_734 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_745(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_742(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_745 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_742 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_750(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_753 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_750 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_761 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_758 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_769 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_766 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_778(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_777 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_774 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_782(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_785 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_782 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_793(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_790(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_793 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_790 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_801(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_798(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_802(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_801 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_798 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_809(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_806(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_809 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_806 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_817(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_814(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_817 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_814 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_825(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_822(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_826(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_825 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_822 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_833(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_830(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_833 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_830 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_841(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_838(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_842(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_841 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_838 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_849(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_846(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_850(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_849 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_846 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_857(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_854(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_858(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_857 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_854 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_865(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_862(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_866(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_865 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_862 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_873(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_870(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_874(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_873 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_870 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_881(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_878(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_882(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_881 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_878 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_889(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_886(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_890(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_889 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_886 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_897(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_894(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_898(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_897 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_894 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_905(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_902(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_906(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_905 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_902 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_913(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_910(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_914(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_913 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_910 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_921(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_918(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_922(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_921 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_918 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_929(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_926(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_930(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_929 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_926 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_937(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_934(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_938(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_937 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_934 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_945(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_942(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_946(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_945 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_942 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_953(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_950(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_954(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_953 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_950 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_961(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_958(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_962(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_961 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_958 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_969(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_966(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_970(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_969 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_966 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_977(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_974(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_978(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_977 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_974 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_985(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_982(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_986(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_985 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_982 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_993(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_990(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_994(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_993 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_990 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_1001(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_998(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_1002(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_1001 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_998 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_1009(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_1006(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_1010(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_1009 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_1006 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_1017(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__2_1014(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__2_1018(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__2_1017 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__2_1014 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__2_2(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__0_116(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__0_117(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__2_2 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__0_116 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__0_118(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__2_50 genblk1_3_a (.a(x[3]), .b(y[3]), .cin(), .sum(s[3]), .carry(
      c1[3]));
   fulladder__2_58 genblk1_4_a (.a(x[4]), .b(y[4]), .cin(), .sum(s1[4]), 
      .carry(c1[4]));
   fulladder__2_66 genblk1_5_a (.a(x[5]), .b(y[5]), .cin(), .sum(s1[5]), 
      .carry(c1[5]));
   fulladder__2_74 genblk1_6_a (.a(x[6]), .b(y[6]), .cin(z[6]), .sum(s1[6]), 
      .carry(c1[6]));
   fulladder__2_82 genblk1_7_a (.a(x[7]), .b(y[7]), .cin(z[7]), .sum(s1[7]), 
      .carry(c1[7]));
   fulladder__2_90 genblk1_8_a (.a(x[8]), .b(y[8]), .cin(z[8]), .sum(s1[8]), 
      .carry(c1[8]));
   fulladder__2_98 genblk1_9_a (.a(x[9]), .b(y[9]), .cin(z[9]), .sum(s1[9]), 
      .carry(c1[9]));
   fulladder__2_106 genblk1_10_a (.a(x[10]), .b(y[10]), .cin(z[10]), .sum(s1[10]), 
      .carry(c1[10]));
   fulladder__2_114 genblk1_11_a (.a(x[11]), .b(y[11]), .cin(z[11]), .sum(s1[11]), 
      .carry(c1[11]));
   fulladder__2_122 genblk1_12_a (.a(x[12]), .b(y[12]), .cin(z[12]), .sum(s1[12]), 
      .carry(c1[12]));
   fulladder__2_130 genblk1_13_a (.a(x[13]), .b(y[13]), .cin(z[13]), .sum(s1[13]), 
      .carry(c1[13]));
   fulladder__2_138 genblk1_14_a (.a(x[14]), .b(y[14]), .cin(z[14]), .sum(s1[14]), 
      .carry(c1[14]));
   fulladder__2_146 genblk1_15_a (.a(x[15]), .b(y[15]), .cin(z[15]), .sum(s1[15]), 
      .carry(c1[15]));
   fulladder__2_154 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(z[16]), .sum(s1[16]), 
      .carry(c1[16]));
   fulladder__2_162 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(z[17]), .sum(s1[17]), 
      .carry(c1[17]));
   fulladder__2_170 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(s1[18]), 
      .carry(c1[18]));
   fulladder__2_178 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(s1[19]), 
      .carry(c1[19]));
   fulladder__2_186 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(s1[20]), 
      .carry(c1[20]));
   fulladder__2_194 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(s1[21]), 
      .carry(c1[21]));
   fulladder__2_202 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(s1[22]), 
      .carry(c1[22]));
   fulladder__2_210 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(s1[23]), 
      .carry(c1[23]));
   fulladder__2_218 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(s1[24]), 
      .carry(c1[24]));
   fulladder__2_226 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(s1[25]), 
      .carry(c1[25]));
   fulladder__2_234 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(s1[26]), 
      .carry(c1[26]));
   fulladder__2_242 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(s1[27]), 
      .carry(c1[27]));
   fulladder__2_250 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(s1[28]), 
      .carry(c1[28]));
   fulladder__2_258 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(s1[29]), 
      .carry(c1[29]));
   fulladder__2_266 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(s1[30]), 
      .carry(c1[30]));
   fulladder__2_274 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(s1[31]), 
      .carry(c1[31]));
   fulladder__2_282 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(s1[32]), 
      .carry(c1[32]));
   fulladder__2_290 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(s1[33]), 
      .carry(c1[33]));
   fulladder__2_298 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(s1[34]), 
      .carry(c1[34]));
   fulladder__2_306 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(s1[35]), 
      .carry(c1[35]));
   fulladder__2_314 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(s1[36]), 
      .carry(c1[36]));
   fulladder__2_322 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(s1[37]), 
      .carry(c1[37]));
   fulladder__2_330 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(s1[38]), 
      .carry(c1[38]));
   fulladder__2_338 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(s1[39]), 
      .carry(c1[39]));
   fulladder__2_346 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(s1[40]), 
      .carry(c1[40]));
   fulladder__2_354 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(s1[41]), 
      .carry(c1[41]));
   fulladder__2_362 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(s1[42]), 
      .carry(c1[42]));
   fulladder__2_370 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(s1[43]), 
      .carry(c1[43]));
   fulladder__2_378 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(s1[44]), 
      .carry(c1[44]));
   fulladder__2_386 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(s1[45]), 
      .carry(c1[45]));
   fulladder__2_394 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(s1[46]), 
      .carry(c1[46]));
   fulladder__2_402 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(s1[47]), 
      .carry(c1[47]));
   fulladder__2_410 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(s1[48]), 
      .carry(c1[48]));
   fulladder__2_418 genblk1_49_a (.a(x[49]), .b(y[49]), .cin(z[49]), .sum(s1[49]), 
      .carry(c1[49]));
   fulladder__2_426 genblk1_50_a (.a(x[50]), .b(y[50]), .cin(z[50]), .sum(s1[50]), 
      .carry(c1[50]));
   fulladder__2_434 genblk1_51_a (.a(x[51]), .b(y[51]), .cin(z[51]), .sum(s1[51]), 
      .carry(c1[51]));
   fulladder__2_442 genblk1_52_a (.a(x[52]), .b(y[52]), .cin(z[52]), .sum(s1[52]), 
      .carry(c1[52]));
   fulladder__2_450 genblk1_53_a (.a(x[53]), .b(y[53]), .cin(z[53]), .sum(s1[53]), 
      .carry(c1[53]));
   fulladder__2_458 genblk1_54_a (.a(x[54]), .b(y[54]), .cin(z[54]), .sum(s1[54]), 
      .carry(c1[54]));
   fulladder__2_466 genblk1_55_a (.a(x[55]), .b(y[55]), .cin(z[55]), .sum(s1[55]), 
      .carry(c1[55]));
   fulladder__2_474 genblk1_56_a (.a(x[56]), .b(y[56]), .cin(z[56]), .sum(s1[56]), 
      .carry(c1[56]));
   fulladder__2_482 genblk1_57_a (.a(x[57]), .b(y[57]), .cin(z[57]), .sum(s1[57]), 
      .carry(c1[57]));
   fulladder__2_490 genblk1_58_a (.a(x[58]), .b(y[58]), .cin(z[58]), .sum(s1[58]), 
      .carry(c1[58]));
   fulladder__2_498 genblk1_59_a (.a(x[59]), .b(y[59]), .cin(z[59]), .sum(s1[59]), 
      .carry(c1[59]));
   fulladder__2_506 genblk1_60_a (.a(x[60]), .b(y[60]), .cin(z[60]), .sum(s1[60]), 
      .carry(c1[60]));
   fulladder__2_514 genblk1_61_a (.a(x[61]), .b(y[61]), .cin(z[61]), .sum(s1[61]), 
      .carry(c1[61]));
   fulladder__2_522 genblk1_62_a (.a(x[62]), .b(y[62]), .cin(z[62]), .sum(s1[62]), 
      .carry(c1[62]));
   fulladder__2_530 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[63]), 
      .carry());
   fulladder__2_554 genblk2_3_b (.a(s1[4]), .b(c1[3]), .cin(), .sum(s[4]), 
      .carry(c2[4]));
   fulladder__2_562 genblk2_4_b (.a(s1[5]), .b(c1[4]), .cin(c2[4]), .sum(s[5]), 
      .carry(c2[5]));
   fulladder__2_570 genblk2_5_b (.a(s1[6]), .b(c1[5]), .cin(c2[5]), .sum(s[6]), 
      .carry(c2[6]));
   fulladder__2_578 genblk2_6_b (.a(s1[7]), .b(c1[6]), .cin(c2[6]), .sum(s[7]), 
      .carry(c2[7]));
   fulladder__2_586 genblk2_7_b (.a(s1[8]), .b(c1[7]), .cin(c2[7]), .sum(s[8]), 
      .carry(c2[8]));
   fulladder__2_594 genblk2_8_b (.a(s1[9]), .b(c1[8]), .cin(c2[8]), .sum(s[9]), 
      .carry(c2[9]));
   fulladder__2_602 genblk2_9_b (.a(s1[10]), .b(c1[9]), .cin(c2[9]), .sum(s[10]), 
      .carry(c2[10]));
   fulladder__2_610 genblk2_10_b (.a(s1[11]), .b(c1[10]), .cin(c2[10]), .sum(
      s[11]), .carry(c2[11]));
   fulladder__2_618 genblk2_11_b (.a(s1[12]), .b(c1[11]), .cin(c2[11]), .sum(
      s[12]), .carry(c2[12]));
   fulladder__2_626 genblk2_12_b (.a(s1[13]), .b(c1[12]), .cin(c2[12]), .sum(
      s[13]), .carry(c2[13]));
   fulladder__2_634 genblk2_13_b (.a(s1[14]), .b(c1[13]), .cin(c2[13]), .sum(
      s[14]), .carry(c2[14]));
   fulladder__2_642 genblk2_14_b (.a(s1[15]), .b(c1[14]), .cin(c2[14]), .sum(
      s[15]), .carry(c2[15]));
   fulladder__2_650 genblk2_15_b (.a(s1[16]), .b(c1[15]), .cin(c2[15]), .sum(
      s[16]), .carry(c2[16]));
   fulladder__2_658 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(c2[16]), .sum(
      s[17]), .carry(c2[17]));
   fulladder__2_666 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), .sum(
      s[18]), .carry(c2[18]));
   fulladder__2_674 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), .sum(
      s[19]), .carry(c2[19]));
   fulladder__2_682 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), .sum(
      s[20]), .carry(c2[20]));
   fulladder__2_690 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), .sum(
      s[21]), .carry(c2[21]));
   fulladder__2_698 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), .sum(
      s[22]), .carry(c2[22]));
   fulladder__2_706 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), .sum(
      s[23]), .carry(c2[23]));
   fulladder__2_714 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), .sum(
      s[24]), .carry(c2[24]));
   fulladder__2_722 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), .sum(
      s[25]), .carry(c2[25]));
   fulladder__2_730 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), .sum(
      s[26]), .carry(c2[26]));
   fulladder__2_738 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), .sum(
      s[27]), .carry(c2[27]));
   fulladder__2_746 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), .sum(
      s[28]), .carry(c2[28]));
   fulladder__2_754 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), .sum(
      s[29]), .carry(c2[29]));
   fulladder__2_762 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), .sum(
      s[30]), .carry(c2[30]));
   fulladder__2_770 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), .sum(
      s[31]), .carry(c2[31]));
   fulladder__2_778 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), .sum(
      s[32]), .carry(c2[32]));
   fulladder__2_786 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), .sum(
      s[33]), .carry(c2[33]));
   fulladder__2_794 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), .sum(
      s[34]), .carry(c2[34]));
   fulladder__2_802 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), .sum(
      s[35]), .carry(c2[35]));
   fulladder__2_810 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), .sum(
      s[36]), .carry(c2[36]));
   fulladder__2_818 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), .sum(
      s[37]), .carry(c2[37]));
   fulladder__2_826 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), .sum(
      s[38]), .carry(c2[38]));
   fulladder__2_834 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), .sum(
      s[39]), .carry(c2[39]));
   fulladder__2_842 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), .sum(
      s[40]), .carry(c2[40]));
   fulladder__2_850 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), .sum(
      s[41]), .carry(c2[41]));
   fulladder__2_858 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), .sum(
      s[42]), .carry(c2[42]));
   fulladder__2_866 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), .sum(
      s[43]), .carry(c2[43]));
   fulladder__2_874 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), .sum(
      s[44]), .carry(c2[44]));
   fulladder__2_882 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), .sum(
      s[45]), .carry(c2[45]));
   fulladder__2_890 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), .sum(
      s[46]), .carry(c2[46]));
   fulladder__2_898 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), .sum(
      s[47]), .carry(c2[47]));
   fulladder__2_906 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), .sum(
      s[48]), .carry(c2[48]));
   fulladder__2_914 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), .sum(
      s[49]), .carry(c2[49]));
   fulladder__2_922 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), .sum(
      s[50]), .carry(c2[50]));
   fulladder__2_930 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), .sum(
      s[51]), .carry(c2[51]));
   fulladder__2_938 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), .sum(
      s[52]), .carry(c2[52]));
   fulladder__2_946 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), .sum(
      s[53]), .carry(c2[53]));
   fulladder__2_954 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), .sum(
      s[54]), .carry(c2[54]));
   fulladder__2_962 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), .sum(
      s[55]), .carry(c2[55]));
   fulladder__2_970 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), .sum(
      s[56]), .carry(c2[56]));
   fulladder__2_978 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), .sum(
      s[57]), .carry(c2[57]));
   fulladder__2_986 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), .sum(
      s[58]), .carry(c2[58]));
   fulladder__2_994 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), .sum(
      s[59]), .carry(c2[59]));
   fulladder__2_1002 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__2_1010 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__2_1018 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__0_117 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), .sum(
      s[63]), .carry());
endmodule

module halfadder__3_225(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_226(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__3_225 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__3_233(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_230(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_234(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_233 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_230 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_241(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_238(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_241 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_238 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_246(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_249 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_246 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_258(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_257 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_254 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_265 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_262 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_273 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_270 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_278(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_281 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_278 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_289(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_286(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_289 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_286 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_297(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_294(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_298(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_297 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_294 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_305(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_302(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_306(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_305 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_302 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_313(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_310(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_313 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_310 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_321(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_318(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_322(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_321 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_318 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_329(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_326(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_330(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_329 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_326 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_337(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_334(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_337 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_334 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_345(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_342(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_346(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_345 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_342 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_353(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_350(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_354(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_353 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_350 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_361(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_358(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_362(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_361 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_358 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_369(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_366(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_370(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_369 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_366 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_377(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_374(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_378(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_377 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_374 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_385(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_382(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_386(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_385 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_382 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_393(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_390(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_394(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_393 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_390 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_401(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_398(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_402(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_401 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_398 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_409(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_406(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_410(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_409 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_406 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_417(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_414(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_418(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_417 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_414 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_425(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_422(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_426(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_425 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_422 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_433(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_430(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_434(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_433 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_430 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_441(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_438(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_442(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_441 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_438 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_449(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_446(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_450(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_449 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_446 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_457(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_454(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_458(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_457 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_454 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_465(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_462(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_466(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_465 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_462 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_473(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_470(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_474(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_473 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_470 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_481(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_478(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_482(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_481 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_478 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_489(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_486(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_490(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_489 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_486 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_497(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_494(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_498(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_497 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_494 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_505(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_502(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_506(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_505 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_502 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_513(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_510(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_514(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_513 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_510 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_521 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_518 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__3_526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__3_530(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__3_529 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__3_526 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__3_729(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_730(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__3_729 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__3_737(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_734(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_737 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_734 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_745(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_742(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_745 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_742 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_750(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_753 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_750 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_761 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_758 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_769 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_766 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_778(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_777 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_774 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_782(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_785 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_782 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_793(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_790(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_793 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_790 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_801(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_798(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_802(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_801 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_798 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_809(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_806(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_809 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_806 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_817(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_814(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_817 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_814 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_825(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_822(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_826(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_825 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_822 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_833(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_830(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_833 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_830 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_841(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_838(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_842(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_841 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_838 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_849(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_846(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_850(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_849 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_846 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_857(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_854(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_858(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_857 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_854 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_865(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_862(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_866(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_865 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_862 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_873(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_870(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_874(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_873 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_870 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_881(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_878(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_882(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_881 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_878 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_889(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_886(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_890(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_889 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_886 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_897(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_894(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_898(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_897 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_894 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_905(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_902(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_906(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_905 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_902 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_913(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_910(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_914(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_913 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_910 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_921(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_918(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_922(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_921 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_918 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_929(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_926(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_930(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_929 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_926 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_937(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_934(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_938(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_937 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_934 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_945(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_942(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_946(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_945 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_942 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_953(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_950(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_954(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_953 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_950 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_961(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_958(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_962(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_961 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_958 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_969(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_966(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_970(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_969 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_966 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_977(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_974(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_978(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_977 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_974 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_985(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_982(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_986(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_985 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_982 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_993(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_990(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_994(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_993 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_990 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_1001(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_998(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_1002(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_1001 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_998 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_1009(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_1006(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_1010(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_1009 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_1006 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_1017(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__3_1014(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__3_1018(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__3_1017 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__3_1014 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__3_2(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__0_123(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__0_124(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__3_2 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__0_123 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__0_125(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__3_226 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(), .sum(s[25]), 
      .carry(c1[25]));
   fulladder__3_234 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(s1[26]), 
      .carry(c1[26]));
   fulladder__3_242 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(s1[27]), 
      .carry(c1[27]));
   fulladder__3_250 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(s1[28]), 
      .carry(c1[28]));
   fulladder__3_258 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(s1[29]), 
      .carry(c1[29]));
   fulladder__3_266 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(s1[30]), 
      .carry(c1[30]));
   fulladder__3_274 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(s1[31]), 
      .carry(c1[31]));
   fulladder__3_282 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(s1[32]), 
      .carry(c1[32]));
   fulladder__3_290 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(s1[33]), 
      .carry(c1[33]));
   fulladder__3_298 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(s1[34]), 
      .carry(c1[34]));
   fulladder__3_306 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(s1[35]), 
      .carry(c1[35]));
   fulladder__3_314 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(s1[36]), 
      .carry(c1[36]));
   fulladder__3_322 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(s1[37]), 
      .carry(c1[37]));
   fulladder__3_330 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(s1[38]), 
      .carry(c1[38]));
   fulladder__3_338 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(s1[39]), 
      .carry(c1[39]));
   fulladder__3_346 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(s1[40]), 
      .carry(c1[40]));
   fulladder__3_354 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(s1[41]), 
      .carry(c1[41]));
   fulladder__3_362 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(s1[42]), 
      .carry(c1[42]));
   fulladder__3_370 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(s1[43]), 
      .carry(c1[43]));
   fulladder__3_378 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(s1[44]), 
      .carry(c1[44]));
   fulladder__3_386 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(s1[45]), 
      .carry(c1[45]));
   fulladder__3_394 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(s1[46]), 
      .carry(c1[46]));
   fulladder__3_402 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(s1[47]), 
      .carry(c1[47]));
   fulladder__3_410 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(s1[48]), 
      .carry(c1[48]));
   fulladder__3_418 genblk1_49_a (.a(x[49]), .b(y[49]), .cin(z[49]), .sum(s1[49]), 
      .carry(c1[49]));
   fulladder__3_426 genblk1_50_a (.a(x[50]), .b(y[50]), .cin(z[50]), .sum(s1[50]), 
      .carry(c1[50]));
   fulladder__3_434 genblk1_51_a (.a(x[51]), .b(y[51]), .cin(z[51]), .sum(s1[51]), 
      .carry(c1[51]));
   fulladder__3_442 genblk1_52_a (.a(x[52]), .b(y[52]), .cin(z[52]), .sum(s1[52]), 
      .carry(c1[52]));
   fulladder__3_450 genblk1_53_a (.a(x[53]), .b(y[53]), .cin(z[53]), .sum(s1[53]), 
      .carry(c1[53]));
   fulladder__3_458 genblk1_54_a (.a(x[54]), .b(y[54]), .cin(z[54]), .sum(s1[54]), 
      .carry(c1[54]));
   fulladder__3_466 genblk1_55_a (.a(x[63]), .b(y[55]), .cin(z[55]), .sum(s1[55]), 
      .carry(c1[55]));
   fulladder__3_474 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[56]), .sum(s1[56]), 
      .carry(c1[56]));
   fulladder__3_482 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[57]), 
      .carry(c1[57]));
   fulladder__3_490 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[58]), 
      .carry(c1[58]));
   fulladder__3_498 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[59]), 
      .carry(c1[59]));
   fulladder__3_506 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[60]), 
      .carry(c1[60]));
   fulladder__3_514 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[61]), 
      .carry(c1[61]));
   fulladder__3_522 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[62]), 
      .carry(c1[62]));
   fulladder__3_530 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[63]), 
      .carry());
   fulladder__3_730 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(), .sum(s[26]), 
      .carry(c2[26]));
   fulladder__3_738 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), .sum(
      s[27]), .carry(c2[27]));
   fulladder__3_746 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), .sum(
      s[28]), .carry(c2[28]));
   fulladder__3_754 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), .sum(
      s[29]), .carry(c2[29]));
   fulladder__3_762 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), .sum(
      s[30]), .carry(c2[30]));
   fulladder__3_770 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), .sum(
      s[31]), .carry(c2[31]));
   fulladder__3_778 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), .sum(
      s[32]), .carry(c2[32]));
   fulladder__3_786 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), .sum(
      s[33]), .carry(c2[33]));
   fulladder__3_794 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), .sum(
      s[34]), .carry(c2[34]));
   fulladder__3_802 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), .sum(
      s[35]), .carry(c2[35]));
   fulladder__3_810 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), .sum(
      s[36]), .carry(c2[36]));
   fulladder__3_818 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), .sum(
      s[37]), .carry(c2[37]));
   fulladder__3_826 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), .sum(
      s[38]), .carry(c2[38]));
   fulladder__3_834 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), .sum(
      s[39]), .carry(c2[39]));
   fulladder__3_842 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), .sum(
      s[40]), .carry(c2[40]));
   fulladder__3_850 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), .sum(
      s[41]), .carry(c2[41]));
   fulladder__3_858 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), .sum(
      s[42]), .carry(c2[42]));
   fulladder__3_866 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), .sum(
      s[43]), .carry(c2[43]));
   fulladder__3_874 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), .sum(
      s[44]), .carry(c2[44]));
   fulladder__3_882 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), .sum(
      s[45]), .carry(c2[45]));
   fulladder__3_890 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), .sum(
      s[46]), .carry(c2[46]));
   fulladder__3_898 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), .sum(
      s[47]), .carry(c2[47]));
   fulladder__3_906 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), .sum(
      s[48]), .carry(c2[48]));
   fulladder__3_914 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), .sum(
      s[49]), .carry(c2[49]));
   fulladder__3_922 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), .sum(
      s[50]), .carry(c2[50]));
   fulladder__3_930 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), .sum(
      s[51]), .carry(c2[51]));
   fulladder__3_938 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), .sum(
      s[52]), .carry(c2[52]));
   fulladder__3_946 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), .sum(
      s[53]), .carry(c2[53]));
   fulladder__3_954 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), .sum(
      s[54]), .carry(c2[54]));
   fulladder__3_962 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), .sum(
      s[55]), .carry(c2[55]));
   fulladder__3_970 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), .sum(
      s[56]), .carry(c2[56]));
   fulladder__3_978 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), .sum(
      s[57]), .carry(c2[57]));
   fulladder__3_986 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), .sum(
      s[58]), .carry(c2[58]));
   fulladder__3_994 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), .sum(
      s[59]), .carry(c2[59]));
   fulladder__3_1002 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__3_1010 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__3_1018 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__0_124 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), .sum(
      s[63]), .carry());
endmodule

module halfadder__4_1849(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1850(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_1849 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_1841(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1838(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1842(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1841 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1838 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1833(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1830(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1833 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1830 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1825(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1822(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1826(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1825 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1822 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1817(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1814(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1817 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1814 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1809(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1806(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1809 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1806 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1801(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1798(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1802(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1801 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1798 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1793(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1790(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1793 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1790 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1782(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1785 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1782 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1778(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1777 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1774 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1769 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1766 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1761 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1758 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1750(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1753 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1750 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1745(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1742(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1745 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1742 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1737(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1734(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1737 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1734 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1729(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1726(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1730(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1729 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1726 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1721(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1718(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1722(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1721 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1718 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1713(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1710(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1714(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1713 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1710 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1705(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1702(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1706(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1705 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1702 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1697(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1694(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1698(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1697 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1694 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1689(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1686(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1690(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1689 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1686 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1681(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1678(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1682(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1681 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1678 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1673(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1670(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1674(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1673 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1670 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1665(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1662(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1666(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1665 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1662 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1657(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1654(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1658(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1657 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1654 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1649(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1646(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1650(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1649 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1646 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1641(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1638(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1642(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1641 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1638 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1633(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1630(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1634(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1633 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1630 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1625(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1622(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1626(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1625 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1622 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1617(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1614(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1618(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1617 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1614 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1609(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1606(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1610(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1609 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1606 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1601(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1598(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1602(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1601 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1598 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1593(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1590(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1594(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1593 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1590 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1585(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1582(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1586(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1585 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1582 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1577(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1574(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1578(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1577 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1574 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1569(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1566(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1570(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1569 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1566 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1561(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1558(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1562(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1561 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1558 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1553(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1550(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1554(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1553 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1550 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1545(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1542(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1546(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1545 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1542 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1537(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1534(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1538(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1537 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1534 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1530(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1529 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1526 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__4_1518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__4_1522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__4_1521 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__4_1518 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__4_1345(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1346(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_1345 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_1337(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1334(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1337 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1334 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1329(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1326(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1330(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1329 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1326 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1321(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1318(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1322(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1321 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1318 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1313(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1310(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1313 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1310 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1305(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1302(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1306(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1305 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1302 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1297(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1294(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1298(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1297 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1294 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1289(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1286(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1289 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1286 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1278(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1281 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1278 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1273 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1270 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1265 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1262 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1258(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1257 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1254 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1246(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1249 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1246 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1241(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1238(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1241 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1238 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1233(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1230(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1234(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1233 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1230 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1225(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1222(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1226(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1225 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1222 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1217(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1214(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1217 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1214 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1209(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1206(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1210(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1209 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1206 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1201(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1198(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1202(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1201 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1198 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1193(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1190(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1194(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1193 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1190 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1185(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1182(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1186(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1185 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1182 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1177(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1174(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1178(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1177 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1174 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1169(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1166(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1170(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1169 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1166 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1161(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1158(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1162(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1161 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1158 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1153(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1150(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1154(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1153 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1150 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1145(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1142(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1146(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1145 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1142 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1137(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1134(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1138(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1137 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1134 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1129(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1126(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1130(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1129 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1126 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1121(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1118(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1122(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1121 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1118 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1113(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1110(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1114(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1113 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1110 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1105(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1102(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1106(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1105 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1102 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1097(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1094(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1098(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1097 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1094 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1089(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1086(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1090(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1089 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1086 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1081(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1078(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1082(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1081 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1078 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1073(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1070(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1074(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1073 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1070 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1065(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1062(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1066(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1065 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1062 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1057(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1054(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1058(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1057 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1054 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1049(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1046(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1050(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1049 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1046 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1041(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1038(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1042(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1041 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1038 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1033(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1030(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1034(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1033 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1030 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1025(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__4_1022(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__4_1026(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__4_1025 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__4_1022 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__4_2043(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__4_1850 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(), .sum(s[22]), 
      .carry(c1[22]));
   fulladder__4_1842 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__4_1834 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__4_1826 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__4_1818 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__4_1810 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__4_1802 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__4_1794 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__4_1786 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__4_1778 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__4_1770 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__4_1762 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__4_1754 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__4_1746 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__4_1738 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__4_1730 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__4_1722 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__4_1714 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__4_1706 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__4_1698 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__4_1690 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__4_1682 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__4_1674 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__4_1666 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__4_1658 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__4_1650 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__4_1642 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__4_1634 genblk1_49_a (.a(x[49]), .b(y[49]), .cin(z[49]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__4_1626 genblk1_50_a (.a(x[50]), .b(y[50]), .cin(z[50]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__4_1618 genblk1_51_a (.a(x[51]), .b(y[51]), .cin(z[51]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__4_1610 genblk1_52_a (.a(x[63]), .b(y[52]), .cin(z[52]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__4_1602 genblk1_53_a (.a(x[63]), .b(y[63]), .cin(z[53]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__4_1594 genblk1_54_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__4_1586 genblk1_55_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__4_1578 genblk1_56_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__4_1570 genblk1_57_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__4_1562 genblk1_58_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__4_1554 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__4_1546 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__4_1538 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__4_1530 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__4_1522 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__4_1346 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(), .sum(s[23]), 
      .carry(c2[23]));
   fulladder__4_1338 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__4_1330 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__4_1322 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__4_1314 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__4_1306 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__4_1298 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__4_1290 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__4_1282 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__4_1274 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__4_1266 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__4_1258 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__4_1250 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__4_1242 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__4_1234 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__4_1226 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__4_1218 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__4_1210 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__4_1202 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__4_1194 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__4_1186 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__4_1178 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__4_1170 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__4_1162 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__4_1154 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__4_1146 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__4_1138 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__4_1130 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__4_1122 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__4_1114 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__4_1106 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__4_1098 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__4_1090 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__4_1082 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__4_1074 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__4_1066 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__4_1058 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__4_1050 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__4_1042 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__4_1034 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__4_1026 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__4_2978(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2979(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2978 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2970(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2971(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2970 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2962(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2963(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2962 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2954(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2955(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2954 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2946(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2947(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2946 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2938(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2939(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2938 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2930(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2931(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2930 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2922(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2923(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2922 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2914(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2915(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2914 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2906(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2903(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2907(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2906 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2903 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2898(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2895(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2899(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2898 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2895 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2890(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2887(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2891(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2890 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2887 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2882(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2879(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2883(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2882 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2879 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2874(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2871(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2875(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2874 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2871 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2866(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2863(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2867(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2866 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2863 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2858(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2855(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2859(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2858 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2855 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2850(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2847(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2851(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2850 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2847 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2842(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2839(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2843(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2842 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2839 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2834(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2831(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2835(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2834 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2831 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2826(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2823(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2827(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2826 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2823 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2818(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2815(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2819(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2818 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2815 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2810(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2807(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2811(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2810 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2807 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2802(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2799(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2803(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2802 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2799 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2794(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2791(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2795(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2794 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2791 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2786(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2783(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2787(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2786 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2783 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2778(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2775(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2779(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2778 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2775 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2770(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2767(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2771(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2770 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2767 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2762(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2759(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2763(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2762 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2759 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2754(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2751(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2755(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2754 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2751 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2746(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2743(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2747(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2746 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2743 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2738(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2735(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2739(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2738 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2735 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2730(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2727(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2731(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2730 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2727 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2722(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2719(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2723(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2722 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2719 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2714(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2711(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2715(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2714 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2711 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2706(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2703(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2707(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2706 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2703 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2698(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2695(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2699(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2698 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2695 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2690(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2687(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2691(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2690 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2687 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2682(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2679(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2683(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2682 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2679 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2674(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2671(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2675(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2674 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2671 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2666(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2663(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2667(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2666 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2663 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2658(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2655(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2659(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2658 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2655 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2650(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2647(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2651(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2650 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2647 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2642(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2639(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2643(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2642 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2639 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2634(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2631(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2635(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2634 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2631 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2626(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2623(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2627(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2626 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2623 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2618(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2615(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2619(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2618 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2615 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2610(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2607(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2611(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2610 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2607 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2602(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2599(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2603(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2602 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2599 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2594(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2591(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2595(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2594 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2591 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2586(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2583(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2587(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2586 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2583 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2578(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2575(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2579(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2578 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2575 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2570(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2567(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2571(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2570 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2567 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2562(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2559(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2563(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2562 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2559 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2554(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2551(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2555(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2554 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2551 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2546(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__4_2543(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__4_2547(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__4_2546 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__4_2543 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__4_2474(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2475(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_2474 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_2466(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2463(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2467(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2466 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2463 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2458(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2455(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2459(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2458 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2455 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2450(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2447(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2451(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2450 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2447 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2442(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2439(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2443(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2442 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2439 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2434(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2431(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2435(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2434 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2431 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2426(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2423(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2427(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2426 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2423 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2418(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2415(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2419(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2418 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2415 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2410(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2407(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2411(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2410 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2407 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2402(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2399(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2403(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2402 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2399 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2394(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2391(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2395(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2394 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2391 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2386(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2383(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2387(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2386 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2383 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2378(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2375(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2379(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2378 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2375 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2370(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2367(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2371(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2370 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2367 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2362(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2359(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2363(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2362 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2359 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2354(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2351(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2355(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2354 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2351 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2346(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2343(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2347(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2346 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2343 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2338(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2335(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2339(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2338 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2335 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2330(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2327(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2331(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2330 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2327 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2322(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2319(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2323(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2322 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2319 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2314(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2311(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2315(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2314 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2311 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2306(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2303(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2307(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2306 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2303 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2298(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2295(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2299(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2298 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2295 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2290(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2287(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2291(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2290 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2287 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2282(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2279(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2283(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2282 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2279 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2274(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2271(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2275(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2274 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2271 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2266(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2263(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2267(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2266 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2263 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2258(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2255(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2259(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2258 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2255 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2250(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2247(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2251(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2250 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2247 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2242(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2239(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2243(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2242 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2239 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2234(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2231(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2235(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2234 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2231 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2226(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2223(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2227(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2226 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2223 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2218(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2215(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2219(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2218 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2215 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2210(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2207(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2211(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2210 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2207 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2202(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2199(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2203(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2202 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2199 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2194(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2191(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2195(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2194 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2191 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2186(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2183(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2187(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2186 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2183 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2178(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2175(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2179(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2178 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2175 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2170(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2167(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2171(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2170 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2167 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2162(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2159(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2163(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2162 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2159 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2154(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2151(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2155(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2154 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2151 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2146(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2143(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2147(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2146 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2143 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2138(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2135(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2139(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2138 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2135 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2130(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2127(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2131(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2130 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2127 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2122(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2119(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2123(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2122 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2119 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2114(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2111(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2115(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2114 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2111 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2106(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2103(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2107(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2106 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2103 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2098(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2095(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2099(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2098 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2095 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2090(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2087(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2091(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2090 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2087 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2082(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2079(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2083(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2082 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2079 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2074(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2071(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2075(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2074 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2071 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2066(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2063(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2067(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2066 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2063 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2058(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_2055(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_2059(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_2058 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_2055 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2050(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__4_2047(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__4_2051(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__4_2050 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__4_2047 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__4_3068(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__4_2979 genblk1_9_a (.a(x[9]), .b(y[9]), .cin(), .sum(s[9]), 
      .carry(c1[9]));
   fulladder__4_2971 genblk1_10_a (.a(x[10]), .b(y[10]), .cin(), .sum(s1[10]), 
      .carry(c1[10]));
   fulladder__4_2963 genblk1_11_a (.a(x[11]), .b(y[11]), .cin(), .sum(s1[11]), 
      .carry(c1[11]));
   fulladder__4_2955 genblk1_12_a (.a(x[12]), .b(y[12]), .cin(), .sum(s1[12]), 
      .carry(c1[12]));
   fulladder__4_2947 genblk1_13_a (.a(x[13]), .b(y[13]), .cin(), .sum(s1[13]), 
      .carry(c1[13]));
   fulladder__4_2939 genblk1_14_a (.a(x[14]), .b(y[14]), .cin(), .sum(s1[14]), 
      .carry(c1[14]));
   fulladder__4_2931 genblk1_15_a (.a(x[15]), .b(y[15]), .cin(), .sum(s1[15]), 
      .carry(c1[15]));
   fulladder__4_2923 genblk1_16_a (.a(x[16]), .b(y[16]), .cin(), .sum(s1[16]), 
      .carry(c1[16]));
   fulladder__4_2915 genblk1_17_a (.a(x[17]), .b(y[17]), .cin(), .sum(s1[17]), 
      .carry(c1[17]));
   fulladder__4_2907 genblk1_18_a (.a(x[18]), .b(y[18]), .cin(z[18]), .sum(
      s1[18]), .carry(c1[18]));
   fulladder__4_2899 genblk1_19_a (.a(x[19]), .b(y[19]), .cin(z[19]), .sum(
      s1[19]), .carry(c1[19]));
   fulladder__4_2891 genblk1_20_a (.a(x[20]), .b(y[20]), .cin(z[20]), .sum(
      s1[20]), .carry(c1[20]));
   fulladder__4_2883 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(z[21]), .sum(
      s1[21]), .carry(c1[21]));
   fulladder__4_2875 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(z[22]), .sum(
      s1[22]), .carry(c1[22]));
   fulladder__4_2867 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(z[23]), .sum(
      s1[23]), .carry(c1[23]));
   fulladder__4_2859 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(
      s1[24]), .carry(c1[24]));
   fulladder__4_2851 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(
      s1[25]), .carry(c1[25]));
   fulladder__4_2843 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(
      s1[26]), .carry(c1[26]));
   fulladder__4_2835 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(
      s1[27]), .carry(c1[27]));
   fulladder__4_2827 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(
      s1[28]), .carry(c1[28]));
   fulladder__4_2819 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(
      s1[29]), .carry(c1[29]));
   fulladder__4_2811 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(
      s1[30]), .carry(c1[30]));
   fulladder__4_2803 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__4_2795 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__4_2787 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__4_2779 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__4_2771 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__4_2763 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__4_2755 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__4_2747 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__4_2739 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__4_2731 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__4_2723 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__4_2715 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__4_2707 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__4_2699 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__4_2691 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__4_2683 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__4_2675 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__4_2667 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__4_2659 genblk1_49_a (.a(x[49]), .b(y[49]), .cin(z[49]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__4_2651 genblk1_50_a (.a(x[50]), .b(y[50]), .cin(z[50]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__4_2643 genblk1_51_a (.a(x[51]), .b(y[51]), .cin(z[51]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__4_2635 genblk1_52_a (.a(x[52]), .b(y[52]), .cin(z[52]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__4_2627 genblk1_53_a (.a(x[53]), .b(y[53]), .cin(z[53]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__4_2619 genblk1_54_a (.a(x[54]), .b(y[54]), .cin(z[54]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__4_2611 genblk1_55_a (.a(x[55]), .b(y[55]), .cin(z[55]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__4_2603 genblk1_56_a (.a(x[56]), .b(y[56]), .cin(z[56]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__4_2595 genblk1_57_a (.a(x[57]), .b(y[57]), .cin(z[57]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__4_2587 genblk1_58_a (.a(x[58]), .b(y[58]), .cin(z[58]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__4_2579 genblk1_59_a (.a(x[59]), .b(y[59]), .cin(z[59]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__4_2571 genblk1_60_a (.a(x[60]), .b(y[60]), .cin(z[60]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__4_2563 genblk1_61_a (.a(x[61]), .b(y[61]), .cin(z[61]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__4_2555 genblk1_62_a (.a(x[62]), .b(y[62]), .cin(z[62]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__4_2547 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__4_2475 genblk2_9_b (.a(s1[10]), .b(c1[9]), .cin(), .sum(s[10]), 
      .carry(c2[10]));
   fulladder__4_2467 genblk2_10_b (.a(s1[11]), .b(c1[10]), .cin(c2[10]), 
      .sum(s[11]), .carry(c2[11]));
   fulladder__4_2459 genblk2_11_b (.a(s1[12]), .b(c1[11]), .cin(c2[11]), 
      .sum(s[12]), .carry(c2[12]));
   fulladder__4_2451 genblk2_12_b (.a(s1[13]), .b(c1[12]), .cin(c2[12]), 
      .sum(s[13]), .carry(c2[13]));
   fulladder__4_2443 genblk2_13_b (.a(s1[14]), .b(c1[13]), .cin(c2[13]), 
      .sum(s[14]), .carry(c2[14]));
   fulladder__4_2435 genblk2_14_b (.a(s1[15]), .b(c1[14]), .cin(c2[14]), 
      .sum(s[15]), .carry(c2[15]));
   fulladder__4_2427 genblk2_15_b (.a(s1[16]), .b(c1[15]), .cin(c2[15]), 
      .sum(s[16]), .carry(c2[16]));
   fulladder__4_2419 genblk2_16_b (.a(s1[17]), .b(c1[16]), .cin(c2[16]), 
      .sum(s[17]), .carry(c2[17]));
   fulladder__4_2411 genblk2_17_b (.a(s1[18]), .b(c1[17]), .cin(c2[17]), 
      .sum(s[18]), .carry(c2[18]));
   fulladder__4_2403 genblk2_18_b (.a(s1[19]), .b(c1[18]), .cin(c2[18]), 
      .sum(s[19]), .carry(c2[19]));
   fulladder__4_2395 genblk2_19_b (.a(s1[20]), .b(c1[19]), .cin(c2[19]), 
      .sum(s[20]), .carry(c2[20]));
   fulladder__4_2387 genblk2_20_b (.a(s1[21]), .b(c1[20]), .cin(c2[20]), 
      .sum(s[21]), .carry(c2[21]));
   fulladder__4_2379 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(c2[21]), 
      .sum(s[22]), .carry(c2[22]));
   fulladder__4_2371 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), 
      .sum(s[23]), .carry(c2[23]));
   fulladder__4_2363 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), 
      .sum(s[24]), .carry(c2[24]));
   fulladder__4_2355 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), 
      .sum(s[25]), .carry(c2[25]));
   fulladder__4_2347 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), 
      .sum(s[26]), .carry(c2[26]));
   fulladder__4_2339 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), 
      .sum(s[27]), .carry(c2[27]));
   fulladder__4_2331 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), 
      .sum(s[28]), .carry(c2[28]));
   fulladder__4_2323 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), 
      .sum(s[29]), .carry(c2[29]));
   fulladder__4_2315 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), 
      .sum(s[30]), .carry(c2[30]));
   fulladder__4_2307 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), 
      .sum(s[31]), .carry(c2[31]));
   fulladder__4_2299 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__4_2291 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__4_2283 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__4_2275 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__4_2267 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__4_2259 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__4_2251 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__4_2243 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__4_2235 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__4_2227 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__4_2219 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__4_2211 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__4_2203 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__4_2195 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__4_2187 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__4_2179 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__4_2171 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__4_2163 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__4_2155 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__4_2147 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__4_2139 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__4_2131 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__4_2123 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__4_2115 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__4_2107 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__4_2099 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__4_2091 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__4_2083 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__4_2075 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__4_2067 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__4_2059 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__4_2051 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module halfadder__4_193(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_194(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_193 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_201(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_202(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_201 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_209(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_210(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_209 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_217(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_214(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_217 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_214 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_225(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_222(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_226(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_225 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_222 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_233(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_230(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_234(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_233 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_230 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_241(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_238(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_241 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_238 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_246(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_249 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_246 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_258(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_257 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_254 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_265 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_262 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_273 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_270 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_278(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_281 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_278 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_289(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_286(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_289 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_286 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_297(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_294(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_298(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_297 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_294 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_305(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_302(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_306(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_305 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_302 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_313(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_310(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_313 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_310 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_321(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_318(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_322(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_321 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_318 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_329(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_326(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_330(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_329 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_326 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_337(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_334(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_337 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_334 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_345(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_342(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_346(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_345 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_342 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_353(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_350(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_354(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_353 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_350 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_361(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_358(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_362(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_361 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_358 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_369(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_366(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_370(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_369 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_366 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_377(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_374(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_378(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_377 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_374 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_385(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_382(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_386(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_385 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_382 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_393(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_390(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_394(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_393 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_390 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_401(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_398(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_402(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_401 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_398 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_409(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_406(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_410(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_409 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_406 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_417(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_414(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_418(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_417 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_414 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_425(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_422(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_426(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_425 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_422 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_433(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_430(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_434(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_433 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_430 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_441(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_438(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_442(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_441 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_438 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_449(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_446(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_450(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_449 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_446 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_457(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_454(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_458(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_457 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_454 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_465(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_462(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_466(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_465 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_462 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_473(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_470(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_474(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_473 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_470 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_481(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_478(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_482(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_481 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_478 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_489(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_486(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_490(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_489 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_486 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_497(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_494(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_498(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_497 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_494 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_505(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_502(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_506(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_505 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_502 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_513(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_510(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_514(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_513 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_510 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_521 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_518 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__4_526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__4_530(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__4_529 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__4_526 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__4_697(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_698(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__4_697 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__4_705(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_702(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_706(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_705 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_702 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_713(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_710(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_714(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_713 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_710 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_721(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_718(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_722(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_721 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_718 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_729(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_726(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_730(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_729 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_726 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_737(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_734(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_737 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_734 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_745(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_742(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_745 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_742 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_750(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_753 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_750 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_761 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_758 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_769 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_766 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_778(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_777 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_774 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_782(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_785 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_782 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_793(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_790(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_793 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_790 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_801(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_798(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_802(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_801 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_798 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_809(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_806(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_809 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_806 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_817(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_814(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_817 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_814 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_825(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_822(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_826(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_825 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_822 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_833(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_830(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_833 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_830 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_841(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_838(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_842(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_841 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_838 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_849(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_846(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_850(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_849 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_846 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_857(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_854(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_858(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_857 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_854 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_865(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_862(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_866(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_865 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_862 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_873(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_870(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_874(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_873 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_870 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_881(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_878(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_882(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_881 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_878 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_889(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_886(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_890(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_889 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_886 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_897(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_894(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_898(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_897 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_894 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_905(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_902(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_906(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_905 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_902 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_913(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_910(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_914(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_913 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_910 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_921(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_918(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_922(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_921 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_918 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_929(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_926(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_930(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_929 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_926 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_937(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_934(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_938(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_937 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_934 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_945(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_942(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_946(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_945 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_942 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_953(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_950(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_954(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_953 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_950 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_961(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_958(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_962(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_961 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_958 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_969(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_966(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_970(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_969 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_966 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_977(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_974(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_978(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_977 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_974 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_985(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_982(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_986(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_985 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_982 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_993(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_990(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_994(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_993 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_990 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1001(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_998(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1002(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1001 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_998 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1009(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1006(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1010(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1009 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1006 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_1017(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__4_1014(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__4_1018(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__4_1017 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__4_1014 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__4_2(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__0_129(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__0_130(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__4_2 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__0_129 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__0_131(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__4_194 genblk1_21_a (.a(x[21]), .b(y[21]), .cin(), .sum(s[21]), 
      .carry(c1[21]));
   fulladder__4_202 genblk1_22_a (.a(x[22]), .b(y[22]), .cin(), .sum(s1[22]), 
      .carry(c1[22]));
   fulladder__4_210 genblk1_23_a (.a(x[23]), .b(y[23]), .cin(), .sum(s1[23]), 
      .carry(c1[23]));
   fulladder__4_218 genblk1_24_a (.a(x[24]), .b(y[24]), .cin(z[24]), .sum(s1[24]), 
      .carry(c1[24]));
   fulladder__4_226 genblk1_25_a (.a(x[25]), .b(y[25]), .cin(z[25]), .sum(s1[25]), 
      .carry(c1[25]));
   fulladder__4_234 genblk1_26_a (.a(x[26]), .b(y[26]), .cin(z[26]), .sum(s1[26]), 
      .carry(c1[26]));
   fulladder__4_242 genblk1_27_a (.a(x[27]), .b(y[27]), .cin(z[27]), .sum(s1[27]), 
      .carry(c1[27]));
   fulladder__4_250 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(z[28]), .sum(s1[28]), 
      .carry(c1[28]));
   fulladder__4_258 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(s1[29]), 
      .carry(c1[29]));
   fulladder__4_266 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(s1[30]), 
      .carry(c1[30]));
   fulladder__4_274 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(s1[31]), 
      .carry(c1[31]));
   fulladder__4_282 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(s1[32]), 
      .carry(c1[32]));
   fulladder__4_290 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(s1[33]), 
      .carry(c1[33]));
   fulladder__4_298 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(s1[34]), 
      .carry(c1[34]));
   fulladder__4_306 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(s1[35]), 
      .carry(c1[35]));
   fulladder__4_314 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(s1[36]), 
      .carry(c1[36]));
   fulladder__4_322 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(s1[37]), 
      .carry(c1[37]));
   fulladder__4_330 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(s1[38]), 
      .carry(c1[38]));
   fulladder__4_338 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(s1[39]), 
      .carry(c1[39]));
   fulladder__4_346 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(s1[40]), 
      .carry(c1[40]));
   fulladder__4_354 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(s1[41]), 
      .carry(c1[41]));
   fulladder__4_362 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(s1[42]), 
      .carry(c1[42]));
   fulladder__4_370 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(s1[43]), 
      .carry(c1[43]));
   fulladder__4_378 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(s1[44]), 
      .carry(c1[44]));
   fulladder__4_386 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(s1[45]), 
      .carry(c1[45]));
   fulladder__4_394 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(s1[46]), 
      .carry(c1[46]));
   fulladder__4_402 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(s1[47]), 
      .carry(c1[47]));
   fulladder__4_410 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(s1[48]), 
      .carry(c1[48]));
   fulladder__4_418 genblk1_49_a (.a(x[49]), .b(y[49]), .cin(z[49]), .sum(s1[49]), 
      .carry(c1[49]));
   fulladder__4_426 genblk1_50_a (.a(x[50]), .b(y[50]), .cin(z[50]), .sum(s1[50]), 
      .carry(c1[50]));
   fulladder__4_434 genblk1_51_a (.a(x[51]), .b(y[51]), .cin(z[51]), .sum(s1[51]), 
      .carry(c1[51]));
   fulladder__4_442 genblk1_52_a (.a(x[52]), .b(y[52]), .cin(z[52]), .sum(s1[52]), 
      .carry(c1[52]));
   fulladder__4_450 genblk1_53_a (.a(x[53]), .b(y[53]), .cin(z[53]), .sum(s1[53]), 
      .carry(c1[53]));
   fulladder__4_458 genblk1_54_a (.a(x[54]), .b(y[54]), .cin(z[54]), .sum(s1[54]), 
      .carry(c1[54]));
   fulladder__4_466 genblk1_55_a (.a(x[55]), .b(y[55]), .cin(z[55]), .sum(s1[55]), 
      .carry(c1[55]));
   fulladder__4_474 genblk1_56_a (.a(x[56]), .b(y[56]), .cin(z[56]), .sum(s1[56]), 
      .carry(c1[56]));
   fulladder__4_482 genblk1_57_a (.a(x[57]), .b(y[57]), .cin(z[57]), .sum(s1[57]), 
      .carry(c1[57]));
   fulladder__4_490 genblk1_58_a (.a(x[58]), .b(y[58]), .cin(z[58]), .sum(s1[58]), 
      .carry(c1[58]));
   fulladder__4_498 genblk1_59_a (.a(x[59]), .b(y[59]), .cin(z[59]), .sum(s1[59]), 
      .carry(c1[59]));
   fulladder__4_506 genblk1_60_a (.a(x[60]), .b(y[60]), .cin(z[60]), .sum(s1[60]), 
      .carry(c1[60]));
   fulladder__4_514 genblk1_61_a (.a(x[61]), .b(y[61]), .cin(z[61]), .sum(s1[61]), 
      .carry(c1[61]));
   fulladder__4_522 genblk1_62_a (.a(x[62]), .b(y[62]), .cin(z[62]), .sum(s1[62]), 
      .carry(c1[62]));
   fulladder__4_530 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[63]), 
      .carry());
   fulladder__4_698 genblk2_21_b (.a(s1[22]), .b(c1[21]), .cin(), .sum(s[22]), 
      .carry(c2[22]));
   fulladder__4_706 genblk2_22_b (.a(s1[23]), .b(c1[22]), .cin(c2[22]), .sum(
      s[23]), .carry(c2[23]));
   fulladder__4_714 genblk2_23_b (.a(s1[24]), .b(c1[23]), .cin(c2[23]), .sum(
      s[24]), .carry(c2[24]));
   fulladder__4_722 genblk2_24_b (.a(s1[25]), .b(c1[24]), .cin(c2[24]), .sum(
      s[25]), .carry(c2[25]));
   fulladder__4_730 genblk2_25_b (.a(s1[26]), .b(c1[25]), .cin(c2[25]), .sum(
      s[26]), .carry(c2[26]));
   fulladder__4_738 genblk2_26_b (.a(s1[27]), .b(c1[26]), .cin(c2[26]), .sum(
      s[27]), .carry(c2[27]));
   fulladder__4_746 genblk2_27_b (.a(s1[28]), .b(c1[27]), .cin(c2[27]), .sum(
      s[28]), .carry(c2[28]));
   fulladder__4_754 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(c2[28]), .sum(
      s[29]), .carry(c2[29]));
   fulladder__4_762 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), .sum(
      s[30]), .carry(c2[30]));
   fulladder__4_770 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), .sum(
      s[31]), .carry(c2[31]));
   fulladder__4_778 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), .sum(
      s[32]), .carry(c2[32]));
   fulladder__4_786 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), .sum(
      s[33]), .carry(c2[33]));
   fulladder__4_794 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), .sum(
      s[34]), .carry(c2[34]));
   fulladder__4_802 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), .sum(
      s[35]), .carry(c2[35]));
   fulladder__4_810 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), .sum(
      s[36]), .carry(c2[36]));
   fulladder__4_818 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), .sum(
      s[37]), .carry(c2[37]));
   fulladder__4_826 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), .sum(
      s[38]), .carry(c2[38]));
   fulladder__4_834 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), .sum(
      s[39]), .carry(c2[39]));
   fulladder__4_842 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), .sum(
      s[40]), .carry(c2[40]));
   fulladder__4_850 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), .sum(
      s[41]), .carry(c2[41]));
   fulladder__4_858 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), .sum(
      s[42]), .carry(c2[42]));
   fulladder__4_866 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), .sum(
      s[43]), .carry(c2[43]));
   fulladder__4_874 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), .sum(
      s[44]), .carry(c2[44]));
   fulladder__4_882 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), .sum(
      s[45]), .carry(c2[45]));
   fulladder__4_890 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), .sum(
      s[46]), .carry(c2[46]));
   fulladder__4_898 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), .sum(
      s[47]), .carry(c2[47]));
   fulladder__4_906 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), .sum(
      s[48]), .carry(c2[48]));
   fulladder__4_914 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), .sum(
      s[49]), .carry(c2[49]));
   fulladder__4_922 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), .sum(
      s[50]), .carry(c2[50]));
   fulladder__4_930 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), .sum(
      s[51]), .carry(c2[51]));
   fulladder__4_938 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), .sum(
      s[52]), .carry(c2[52]));
   fulladder__4_946 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), .sum(
      s[53]), .carry(c2[53]));
   fulladder__4_954 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), .sum(
      s[54]), .carry(c2[54]));
   fulladder__4_962 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), .sum(
      s[55]), .carry(c2[55]));
   fulladder__4_970 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), .sum(
      s[56]), .carry(c2[56]));
   fulladder__4_978 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), .sum(
      s[57]), .carry(c2[57]));
   fulladder__4_986 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), .sum(
      s[58]), .carry(c2[58]));
   fulladder__4_994 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), .sum(
      s[59]), .carry(c2[59]));
   fulladder__4_1002 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__4_1010 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__4_1018 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__0_130 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), .sum(
      s[63]), .carry());
endmodule

module halfadder__5_1785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__5_1785 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__5_1777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1778(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1777 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1774 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1769 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1766 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1761 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1758 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1750(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1753 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1750 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1745(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1742(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1746(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1745 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1742 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1737(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1734(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1738(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1737 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1734 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1729(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1726(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1730(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1729 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1726 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1721(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1718(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1722(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1721 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1718 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1713(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1710(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1714(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1713 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1710 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1705(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1702(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1706(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1705 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1702 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1697(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1694(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1698(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1697 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1694 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1689(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1686(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1690(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1689 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1686 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1681(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1678(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1682(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1681 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1678 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1673(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1670(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1674(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1673 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1670 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1665(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1662(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1666(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1665 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1662 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1657(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1654(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1658(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1657 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1654 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1649(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1646(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1650(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1649 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1646 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1641(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1638(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1642(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1641 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1638 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1633(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1630(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1634(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1633 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1630 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1625(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1622(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1626(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1625 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1622 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1617(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1614(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1618(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1617 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1614 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1609(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1606(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1610(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1609 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1606 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1601(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1598(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1602(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1601 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1598 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1593(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1590(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1594(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1593 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1590 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1585(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1582(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1586(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1585 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1582 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1577(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1574(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1578(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1577 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1574 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1569(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1566(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1570(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1569 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1566 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1561(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1558(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1562(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1561 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1558 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1553(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1550(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1554(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1553 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1550 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1545(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1542(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1546(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1545 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1542 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1537(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1534(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1538(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1537 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1534 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1530(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1529 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1526 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__5_1518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__5_1522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__5_1521 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__5_1518 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__5_1281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__5_1281 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__5_1273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1273 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1270 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1265 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1262 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1258(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1257 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1254 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1246(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1249 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1246 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1241(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1238(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1242(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1241 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1238 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1233(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1230(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1234(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1233 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1230 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1225(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1222(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1226(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1225 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1222 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1217(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1214(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1218(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1217 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1214 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1209(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1206(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1210(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1209 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1206 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1201(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1198(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1202(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1201 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1198 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1193(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1190(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1194(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1193 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1190 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1185(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1182(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1186(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1185 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1182 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1177(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1174(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1178(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1177 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1174 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1169(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1166(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1170(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1169 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1166 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1161(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1158(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1162(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1161 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1158 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1153(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1150(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1154(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1153 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1150 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1145(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1142(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1146(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1145 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1142 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1137(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1134(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1138(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1137 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1134 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1129(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1126(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1130(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1129 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1126 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1121(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1118(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1122(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1121 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1118 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1113(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1110(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1114(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1113 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1110 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1105(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1102(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1106(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1105 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1102 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1097(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1094(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1098(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1097 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1094 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1089(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1086(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1090(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1089 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1086 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1081(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1078(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1082(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1081 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1078 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1073(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1070(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1074(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1073 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1070 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1065(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1062(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1066(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1065 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1062 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1057(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1054(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1058(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1057 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1054 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1049(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1046(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1050(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1049 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1046 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1041(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1038(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1042(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1041 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1038 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1033(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1030(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1034(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1033 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1030 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1025(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__5_1022(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__5_1026(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__5_1025 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__5_1022 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA__5_2043(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__5_1786 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(), .sum(s[30]), 
      .carry(c1[30]));
   fulladder__5_1778 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(
      s1[31]), .carry(c1[31]));
   fulladder__5_1770 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(
      s1[32]), .carry(c1[32]));
   fulladder__5_1762 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(
      s1[33]), .carry(c1[33]));
   fulladder__5_1754 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(
      s1[34]), .carry(c1[34]));
   fulladder__5_1746 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(
      s1[35]), .carry(c1[35]));
   fulladder__5_1738 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(
      s1[36]), .carry(c1[36]));
   fulladder__5_1730 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(
      s1[37]), .carry(c1[37]));
   fulladder__5_1722 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(
      s1[38]), .carry(c1[38]));
   fulladder__5_1714 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(
      s1[39]), .carry(c1[39]));
   fulladder__5_1706 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(
      s1[40]), .carry(c1[40]));
   fulladder__5_1698 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(
      s1[41]), .carry(c1[41]));
   fulladder__5_1690 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(
      s1[42]), .carry(c1[42]));
   fulladder__5_1682 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(
      s1[43]), .carry(c1[43]));
   fulladder__5_1674 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(
      s1[44]), .carry(c1[44]));
   fulladder__5_1666 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(
      s1[45]), .carry(c1[45]));
   fulladder__5_1658 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(
      s1[46]), .carry(c1[46]));
   fulladder__5_1650 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(
      s1[47]), .carry(c1[47]));
   fulladder__5_1642 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(
      s1[48]), .carry(c1[48]));
   fulladder__5_1634 genblk1_49_a (.a(x[49]), .b(y[49]), .cin(z[49]), .sum(
      s1[49]), .carry(c1[49]));
   fulladder__5_1626 genblk1_50_a (.a(x[50]), .b(y[50]), .cin(z[50]), .sum(
      s1[50]), .carry(c1[50]));
   fulladder__5_1618 genblk1_51_a (.a(x[51]), .b(y[51]), .cin(z[51]), .sum(
      s1[51]), .carry(c1[51]));
   fulladder__5_1610 genblk1_52_a (.a(x[52]), .b(y[52]), .cin(z[52]), .sum(
      s1[52]), .carry(c1[52]));
   fulladder__5_1602 genblk1_53_a (.a(x[53]), .b(y[53]), .cin(z[53]), .sum(
      s1[53]), .carry(c1[53]));
   fulladder__5_1594 genblk1_54_a (.a(x[54]), .b(y[54]), .cin(z[54]), .sum(
      s1[54]), .carry(c1[54]));
   fulladder__5_1586 genblk1_55_a (.a(x[55]), .b(y[55]), .cin(z[55]), .sum(
      s1[55]), .carry(c1[55]));
   fulladder__5_1578 genblk1_56_a (.a(x[56]), .b(y[56]), .cin(z[56]), .sum(
      s1[56]), .carry(c1[56]));
   fulladder__5_1570 genblk1_57_a (.a(x[57]), .b(y[57]), .cin(z[57]), .sum(
      s1[57]), .carry(c1[57]));
   fulladder__5_1562 genblk1_58_a (.a(x[58]), .b(y[58]), .cin(z[58]), .sum(
      s1[58]), .carry(c1[58]));
   fulladder__5_1554 genblk1_59_a (.a(x[59]), .b(y[59]), .cin(z[59]), .sum(
      s1[59]), .carry(c1[59]));
   fulladder__5_1546 genblk1_60_a (.a(x[60]), .b(y[60]), .cin(z[60]), .sum(
      s1[60]), .carry(c1[60]));
   fulladder__5_1538 genblk1_61_a (.a(x[61]), .b(y[63]), .cin(z[61]), .sum(
      s1[61]), .carry(c1[61]));
   fulladder__5_1530 genblk1_62_a (.a(x[62]), .b(y[63]), .cin(z[63]), .sum(
      s1[62]), .carry(c1[62]));
   fulladder__5_1522 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(
      s1[63]), .carry());
   fulladder__5_1282 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(), .sum(s[31]), 
      .carry(c2[31]));
   fulladder__5_1274 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), 
      .sum(s[32]), .carry(c2[32]));
   fulladder__5_1266 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), 
      .sum(s[33]), .carry(c2[33]));
   fulladder__5_1258 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), 
      .sum(s[34]), .carry(c2[34]));
   fulladder__5_1250 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), 
      .sum(s[35]), .carry(c2[35]));
   fulladder__5_1242 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), 
      .sum(s[36]), .carry(c2[36]));
   fulladder__5_1234 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), 
      .sum(s[37]), .carry(c2[37]));
   fulladder__5_1226 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), 
      .sum(s[38]), .carry(c2[38]));
   fulladder__5_1218 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), 
      .sum(s[39]), .carry(c2[39]));
   fulladder__5_1210 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), 
      .sum(s[40]), .carry(c2[40]));
   fulladder__5_1202 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), 
      .sum(s[41]), .carry(c2[41]));
   fulladder__5_1194 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), 
      .sum(s[42]), .carry(c2[42]));
   fulladder__5_1186 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), 
      .sum(s[43]), .carry(c2[43]));
   fulladder__5_1178 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), 
      .sum(s[44]), .carry(c2[44]));
   fulladder__5_1170 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), 
      .sum(s[45]), .carry(c2[45]));
   fulladder__5_1162 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), 
      .sum(s[46]), .carry(c2[46]));
   fulladder__5_1154 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), 
      .sum(s[47]), .carry(c2[47]));
   fulladder__5_1146 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), 
      .sum(s[48]), .carry(c2[48]));
   fulladder__5_1138 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), 
      .sum(s[49]), .carry(c2[49]));
   fulladder__5_1130 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), 
      .sum(s[50]), .carry(c2[50]));
   fulladder__5_1122 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), 
      .sum(s[51]), .carry(c2[51]));
   fulladder__5_1114 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), 
      .sum(s[52]), .carry(c2[52]));
   fulladder__5_1106 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), 
      .sum(s[53]), .carry(c2[53]));
   fulladder__5_1098 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), 
      .sum(s[54]), .carry(c2[54]));
   fulladder__5_1090 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), 
      .sum(s[55]), .carry(c2[55]));
   fulladder__5_1082 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), 
      .sum(s[56]), .carry(c2[56]));
   fulladder__5_1074 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), 
      .sum(s[57]), .carry(c2[57]));
   fulladder__5_1066 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), 
      .sum(s[58]), .carry(c2[58]));
   fulladder__5_1058 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), 
      .sum(s[59]), .carry(c2[59]));
   fulladder__5_1050 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__5_1042 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__5_1034 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder__5_1026 genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), 
      .sum(s[63]), .carry());
endmodule

module full_adder__5_2277(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2273(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2269(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2265(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module ripple_adder__5_2278(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2277 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2273 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2269 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2265 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout());
endmodule

module full_adder__5_2295(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2291(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2287(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2283(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module ripple_adder__5_2296(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2295 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2291 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2287 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2283 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout(cout));
endmodule

module full_adder__5_2313(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2309(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2305(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2301(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module ripple_adder__5_2314(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2313 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2309 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2305 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2301 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout(cout));
endmodule

module full_adder__5_2331(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2327(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2323(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2319(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module ripple_adder__5_2332(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2331 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2327 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2323 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2319 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout(cout));
endmodule

module full_adder__5_2349(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2345(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2341(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2337(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module ripple_adder__5_2350(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2349 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2345 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2341 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2337 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout(cout));
endmodule

module full_adder__5_2367(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2363(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2359(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2355(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module ripple_adder__5_2368(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2367 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2363 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2359 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2355 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout(cout));
endmodule

module full_adder__5_2385(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2381(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2377(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2373(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module ripple_adder__5_2386(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2385 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2381 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2377 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2373 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout(cout));
endmodule

module full_adder__5_2403(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2399(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2395(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2391(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module ripple_adder__5_2404(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2403 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2399 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2395 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2391 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout(cout));
endmodule

module full_adder__5_2421(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module full_adder__5_2417(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2413(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module full_adder__5_2409(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module ripple_adder__5_2422(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2421 genblk1_0_FA (.A(in1[0]), .B(in2[0]), .Cin(), .S(s[0]), 
      .Cout(n_0));
   full_adder__5_2417 genblk1_1_FA (.A(in1[1]), .B(in2[1]), .Cin(n_0), .S(s[1]), 
      .Cout(n_1));
   full_adder__5_2413 genblk1_2_FA (.A(in1[2]), .B(in2[2]), .Cin(n_1), .S(s[2]), 
      .Cout(n_2));
   full_adder__5_2409 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(n_2), .S(s[3]), 
      .Cout(cout));
endmodule

module full_adder__5_2427(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module ripple_adder__5_2440(in1, in2, s, cin, cout, OF);
   input [3:0]in1;
   input [3:0]in2;
   output [3:0]s;
   input cin;
   output cout;
   output OF;

   full_adder__5_2427 genblk1_3_FA (.A(in1[3]), .B(in2[3]), .Cin(), .S(s[3]), 
      .Cout(cout));
endmodule

module half_adder__5_2149(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2146(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2143(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2140(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module incrementor__5_2150(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   wire w;

   half_adder__5_2149 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2146 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2143 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder__5_2140 genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), 
      .c(w));
   OR2_X1 i_0_0 (.A1(cin2), .A2(w), .ZN(cout));
endmodule

module half_adder__5_2163(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2160(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2157(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2154(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module incrementor__5_2164(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   wire w;

   half_adder__5_2163 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2160 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2157 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder__5_2154 genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), 
      .c(w));
   OR2_X1 i_0_0 (.A1(cin2), .A2(w), .ZN(cout));
endmodule

module half_adder__5_2177(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2174(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2171(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2168(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module incrementor__5_2178(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   wire w;

   half_adder__5_2177 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2174 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2171 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder__5_2168 genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), 
      .c(w));
   OR2_X1 i_0_0 (.A1(cin2), .A2(w), .ZN(cout));
endmodule

module half_adder__5_2191(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2188(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2185(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2182(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module incrementor__5_2192(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   wire w;

   half_adder__5_2191 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2188 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2185 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder__5_2182 genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), 
      .c(w));
   OR2_X1 i_0_0 (.A1(cin2), .A2(w), .ZN(cout));
endmodule

module half_adder__5_2205(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2202(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2199(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2196(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module incrementor__5_2206(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   wire w;

   half_adder__5_2205 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2202 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2199 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder__5_2196 genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), 
      .c(w));
   OR2_X1 i_0_0 (.A1(cin2), .A2(w), .ZN(cout));
endmodule

module half_adder__5_2219(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2216(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2213(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2210(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module incrementor__5_2220(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   wire w;

   half_adder__5_2219 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2216 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2213 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder__5_2210 genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), 
      .c(w));
   OR2_X1 i_0_0 (.A1(cin2), .A2(w), .ZN(cout));
endmodule

module half_adder__5_2233(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2230(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2227(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2224(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module incrementor__5_2234(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   wire w;

   half_adder__5_2233 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2230 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2227 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder__5_2224 genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), 
      .c(w));
   OR2_X1 i_0_0 (.A1(cin2), .A2(w), .ZN(cout));
endmodule

module half_adder__5_2247(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2244(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2241(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2238(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module incrementor__5_2248(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   wire w;

   half_adder__5_2247 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2244 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2241 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder__5_2238 genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), 
      .c(w));
   OR2_X1 i_0_0 (.A1(cin2), .A2(w), .ZN(cout));
endmodule

module half_adder__5_2046(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2049(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder__5_2052(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
   AND2_X1 i_0_1 (.A1(in1), .A2(in2), .ZN(c));
endmodule

module half_adder(in1, in2, s, c);
   input in1;
   input in2;
   output s;
   output c;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(s));
endmodule

module incrementor(inS, outS, cin1, cin2, cout);
   input [3:0]inS;
   output [3:0]outS;
   input cin1;
   input cin2;
   output cout;

   half_adder__5_2046 genblk1_0_HA (.in1(inS[0]), .in2(cin1), .s(outS[0]), 
      .c(n_0));
   half_adder__5_2049 genblk1_1_HA (.in1(inS[1]), .in2(n_0), .s(outS[1]), 
      .c(n_1));
   half_adder__5_2052 genblk1_2_HA (.in1(inS[2]), .in2(n_1), .s(outS[2]), 
      .c(n_2));
   half_adder genblk1_3_HA (.in1(inS[3]), .in2(n_2), .s(outS[3]), .c());
endmodule

module carry_increment_adder(in1, in2, s, cin, cout, OF);
   input [63:0]in1;
   input [63:0]in2;
   output [63:0]s;
   input cin;
   output cout;
   output OF;

   ripple_adder__5_2278 genblk1_15_RCA (.in1({in1[63], in1[62], in1[61], in1[60]}), 
      .in2({in2[63], in2[62], in2[61], in2[60]}), .s({n_3, n_2, n_1, n_0}), 
      .cin(), .cout(), .OF());
   ripple_adder__5_2296 genblk1_14_RCA (.in1({in1[59], in1[58], in1[57], in1[56]}), 
      .in2({in2[59], in2[58], in2[57], in2[56]}), .s({n_8, n_7, n_6, n_5}), 
      .cin(), .cout(n_4), .OF());
   ripple_adder__5_2314 genblk1_13_RCA (.in1({in1[55], in1[54], in1[53], in1[52]}), 
      .in2({in2[55], in2[54], in2[53], in2[52]}), .s({n_13, n_12, n_11, n_10}), 
      .cin(), .cout(n_9), .OF());
   ripple_adder__5_2332 genblk1_12_RCA (.in1({in1[51], in1[50], in1[49], in1[48]}), 
      .in2({in2[51], in2[50], in2[49], in2[48]}), .s({n_18, n_17, n_16, n_15}), 
      .cin(), .cout(n_14), .OF());
   ripple_adder__5_2350 genblk1_11_RCA (.in1({in1[47], in1[46], in1[45], in1[44]}), 
      .in2({in2[47], in2[46], in2[45], in2[44]}), .s({n_23, n_22, n_21, n_20}), 
      .cin(), .cout(n_19), .OF());
   ripple_adder__5_2368 genblk1_10_RCA (.in1({in1[43], in1[42], in1[41], in1[40]}), 
      .in2({in2[43], in2[42], in2[41], in2[40]}), .s({n_28, n_27, n_26, n_25}), 
      .cin(), .cout(n_24), .OF());
   ripple_adder__5_2386 genblk1_9_RCA (.in1({in1[39], in1[38], in1[37], in1[36]}), 
      .in2({in2[39], in2[38], in2[37], in2[36]}), .s({n_33, n_32, n_31, n_30}), 
      .cin(), .cout(n_29), .OF());
   ripple_adder__5_2404 genblk1_8_RCA (.in1({in1[35], in1[34], in1[33], in1[32]}), 
      .in2({in2[35], in2[34], in2[33], in2[32]}), .s({n_38, n_37, n_36, n_35}), 
      .cin(), .cout(n_34), .OF());
   ripple_adder__5_2422 genblk1_7_RCA (.in1({in1[31], in1[30], in1[29], in1[28]}), 
      .in2({in2[31], in2[30], in2[29], in2[28]}), .s({n_43, n_42, n_41, n_40}), 
      .cin(), .cout(n_39), .OF());
   ripple_adder__5_2440 genblk1_6_RCA (.in1({in1[27], uc_0, uc_1, uc_2}), 
      .in2({in2[27], uc_3, uc_4, uc_5}), .s({s[27], uc_6, uc_7, uc_8}), .cin(), 
      .cout(n_44), .OF());
   incrementor__5_2150 genblk1_7_inc (.inS({n_43, n_42, n_41, n_40}), .outS({
      s[31], s[30], s[29], s[28]}), .cin1(n_44), .cin2(n_39), .cout(n_45));
   incrementor__5_2164 genblk1_8_inc (.inS({n_38, n_37, n_36, n_35}), .outS({
      s[35], s[34], s[33], s[32]}), .cin1(n_45), .cin2(n_34), .cout(n_46));
   incrementor__5_2178 genblk1_9_inc (.inS({n_33, n_32, n_31, n_30}), .outS({
      s[39], s[38], s[37], s[36]}), .cin1(n_46), .cin2(n_29), .cout(n_47));
   incrementor__5_2192 genblk1_10_inc (.inS({n_28, n_27, n_26, n_25}), .outS({
      s[43], s[42], s[41], s[40]}), .cin1(n_47), .cin2(n_24), .cout(n_48));
   incrementor__5_2206 genblk1_11_inc (.inS({n_23, n_22, n_21, n_20}), .outS({
      s[47], s[46], s[45], s[44]}), .cin1(n_48), .cin2(n_19), .cout(n_49));
   incrementor__5_2220 genblk1_12_inc (.inS({n_18, n_17, n_16, n_15}), .outS({
      s[51], s[50], s[49], s[48]}), .cin1(n_49), .cin2(n_14), .cout(n_50));
   incrementor__5_2234 genblk1_13_inc (.inS({n_13, n_12, n_11, n_10}), .outS({
      s[55], s[54], s[53], s[52]}), .cin1(n_50), .cin2(n_9), .cout(n_51));
   incrementor__5_2248 genblk1_14_inc (.inS({n_8, n_7, n_6, n_5}), .outS({s[59], 
      s[58], s[57], s[56]}), .cin1(n_51), .cin2(n_4), .cout(n_52));
   incrementor genblk1_15_inc (.inS({n_3, n_2, n_1, n_0}), .outS({s[63], s[62], 
      s[61], s[60]}), .cin1(n_52), .cin2(), .cout());
endmodule

module halfadder__5_249(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_250(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__5_249 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__5_257(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_254(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_258(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_257 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_254 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_265(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_262(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_266(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_265 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_262 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_273(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_270(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_274(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_273 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_270 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_281(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_278(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_282(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_281 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_278 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_289(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_286(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_290(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_289 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_286 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_297(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_294(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_298(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_297 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_294 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_305(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_302(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_306(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_305 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_302 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_313(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_310(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_314(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_313 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_310 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_321(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_318(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_322(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_321 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_318 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_329(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_326(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_330(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_329 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_326 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_337(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_334(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_338(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_337 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_334 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_345(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_342(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_346(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_345 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_342 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_353(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_350(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_354(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_353 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_350 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_361(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_358(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_362(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_361 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_358 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_369(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_366(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_370(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_369 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_366 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_377(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_374(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_378(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_377 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_374 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_385(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_382(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_386(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_385 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_382 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_393(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_390(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_394(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_393 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_390 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_401(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_398(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_402(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_401 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_398 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_409(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_406(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_410(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_409 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_406 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_417(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_414(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_418(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_417 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_414 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_425(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_422(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_426(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_425 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_422 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_433(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_430(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_434(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_433 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_430 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_441(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_438(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_442(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_441 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_438 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_449(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_446(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_450(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_449 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_446 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_457(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_454(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_458(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_457 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_454 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_465(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_462(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_466(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_465 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_462 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_473(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_470(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_474(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_473 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_470 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_481(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_478(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_482(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_481 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_478 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_489(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_486(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_490(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_489 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_486 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_497(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_494(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_498(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_497 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_494 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_505(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_502(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_506(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_505 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_502 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_513(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_510(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_514(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_513 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_510 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_521(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_518(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_522(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_521 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_518 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_529(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder__5_526(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder__5_530(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__5_529 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder__5_526 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module halfadder__5_753(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_754(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   halfadder__5_753 ha1 (.a(a), .b(b), .sum(sum), .carry(carry));
endmodule

module halfadder__5_761(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_758(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_762(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_761 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_758 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_769(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_766(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_770(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_769 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_766 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_777(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_774(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_778(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_777 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_774 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_785(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_782(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_786(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_785 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_782 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_793(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_790(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_794(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_793 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_790 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_801(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_798(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_802(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_801 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_798 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_809(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_806(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_810(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_809 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_806 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_817(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_814(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_818(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_817 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_814 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_825(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_822(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_826(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_825 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_822 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_833(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_830(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_834(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_833 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_830 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_841(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_838(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_842(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_841 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_838 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_849(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_846(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_850(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_849 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_846 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_857(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_854(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_858(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_857 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_854 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_865(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_862(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_866(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_865 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_862 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_873(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_870(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_874(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_873 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_870 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_881(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_878(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_882(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_881 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_878 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_889(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_886(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_890(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_889 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_886 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_897(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_894(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_898(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_897 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_894 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_905(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_902(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_906(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_905 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_902 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_913(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_910(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_914(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_913 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_910 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_921(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_918(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_922(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_921 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_918 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_929(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_926(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_930(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_929 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_926 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_937(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_934(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_938(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_937 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_934 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_945(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_942(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_946(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_945 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_942 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_953(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_950(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_954(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_953 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_950 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_961(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_958(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_962(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_961 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_958 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_969(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_966(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_970(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_969 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_966 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_977(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_974(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_978(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_977 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_974 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_985(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_982(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_986(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_985 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_982 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_993(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_990(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_994(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_993 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_990 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1001(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_998(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1002(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1001 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_998 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1009(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1006(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1010(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1009 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1006 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_1017(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module halfadder__5_1014(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
   AND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(carry));
endmodule

module fulladder__5_1018(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_carry1;
   wire ha_sum1;
   wire ha_carry2;

   halfadder__5_1017 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry(ha_carry1));
   halfadder__5_1014 ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry(ha_carry2));
   OR2_X1 i_0_0 (.A1(ha_carry1), .A2(ha_carry2), .ZN(carry));
endmodule

module halfadder__5_2(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module halfadder(a, b, sum, carry);
   input a;
   input b;
   output sum;
   output carry;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(sum));
endmodule

module fulladder(a, b, cin, sum, carry);
   input a;
   input b;
   input cin;
   output sum;
   output carry;

   wire ha_sum1;

   halfadder__5_2 ha1 (.a(a), .b(b), .sum(ha_sum1), .carry());
   halfadder ha2 (.a(cin), .b(ha_sum1), .sum(sum), .carry());
endmodule

module CSA(x, y, z, s, carry_final);
   input [63:0]x;
   input [63:0]y;
   input [63:0]z;
   output [63:0]s;
   output [1:0]carry_final;

   wire [63:0]c1;
   wire [63:0]s1;
   wire [63:0]c2;

   fulladder__5_250 genblk1_28_a (.a(x[28]), .b(y[28]), .cin(), .sum(s[28]), 
      .carry(c1[28]));
   fulladder__5_258 genblk1_29_a (.a(x[29]), .b(y[29]), .cin(z[29]), .sum(s1[29]), 
      .carry(c1[29]));
   fulladder__5_266 genblk1_30_a (.a(x[30]), .b(y[30]), .cin(z[30]), .sum(s1[30]), 
      .carry(c1[30]));
   fulladder__5_274 genblk1_31_a (.a(x[31]), .b(y[31]), .cin(z[31]), .sum(s1[31]), 
      .carry(c1[31]));
   fulladder__5_282 genblk1_32_a (.a(x[32]), .b(y[32]), .cin(z[32]), .sum(s1[32]), 
      .carry(c1[32]));
   fulladder__5_290 genblk1_33_a (.a(x[33]), .b(y[33]), .cin(z[33]), .sum(s1[33]), 
      .carry(c1[33]));
   fulladder__5_298 genblk1_34_a (.a(x[34]), .b(y[34]), .cin(z[34]), .sum(s1[34]), 
      .carry(c1[34]));
   fulladder__5_306 genblk1_35_a (.a(x[35]), .b(y[35]), .cin(z[35]), .sum(s1[35]), 
      .carry(c1[35]));
   fulladder__5_314 genblk1_36_a (.a(x[36]), .b(y[36]), .cin(z[36]), .sum(s1[36]), 
      .carry(c1[36]));
   fulladder__5_322 genblk1_37_a (.a(x[37]), .b(y[37]), .cin(z[37]), .sum(s1[37]), 
      .carry(c1[37]));
   fulladder__5_330 genblk1_38_a (.a(x[38]), .b(y[38]), .cin(z[38]), .sum(s1[38]), 
      .carry(c1[38]));
   fulladder__5_338 genblk1_39_a (.a(x[39]), .b(y[39]), .cin(z[39]), .sum(s1[39]), 
      .carry(c1[39]));
   fulladder__5_346 genblk1_40_a (.a(x[40]), .b(y[40]), .cin(z[40]), .sum(s1[40]), 
      .carry(c1[40]));
   fulladder__5_354 genblk1_41_a (.a(x[41]), .b(y[41]), .cin(z[41]), .sum(s1[41]), 
      .carry(c1[41]));
   fulladder__5_362 genblk1_42_a (.a(x[42]), .b(y[42]), .cin(z[42]), .sum(s1[42]), 
      .carry(c1[42]));
   fulladder__5_370 genblk1_43_a (.a(x[43]), .b(y[43]), .cin(z[43]), .sum(s1[43]), 
      .carry(c1[43]));
   fulladder__5_378 genblk1_44_a (.a(x[44]), .b(y[44]), .cin(z[44]), .sum(s1[44]), 
      .carry(c1[44]));
   fulladder__5_386 genblk1_45_a (.a(x[45]), .b(y[45]), .cin(z[45]), .sum(s1[45]), 
      .carry(c1[45]));
   fulladder__5_394 genblk1_46_a (.a(x[46]), .b(y[46]), .cin(z[46]), .sum(s1[46]), 
      .carry(c1[46]));
   fulladder__5_402 genblk1_47_a (.a(x[47]), .b(y[47]), .cin(z[47]), .sum(s1[47]), 
      .carry(c1[47]));
   fulladder__5_410 genblk1_48_a (.a(x[48]), .b(y[48]), .cin(z[48]), .sum(s1[48]), 
      .carry(c1[48]));
   fulladder__5_418 genblk1_49_a (.a(x[49]), .b(y[49]), .cin(z[49]), .sum(s1[49]), 
      .carry(c1[49]));
   fulladder__5_426 genblk1_50_a (.a(x[50]), .b(y[50]), .cin(z[50]), .sum(s1[50]), 
      .carry(c1[50]));
   fulladder__5_434 genblk1_51_a (.a(x[51]), .b(y[51]), .cin(z[51]), .sum(s1[51]), 
      .carry(c1[51]));
   fulladder__5_442 genblk1_52_a (.a(x[52]), .b(y[52]), .cin(z[52]), .sum(s1[52]), 
      .carry(c1[52]));
   fulladder__5_450 genblk1_53_a (.a(x[53]), .b(y[53]), .cin(z[53]), .sum(s1[53]), 
      .carry(c1[53]));
   fulladder__5_458 genblk1_54_a (.a(x[54]), .b(y[54]), .cin(z[54]), .sum(s1[54]), 
      .carry(c1[54]));
   fulladder__5_466 genblk1_55_a (.a(x[55]), .b(y[55]), .cin(z[55]), .sum(s1[55]), 
      .carry(c1[55]));
   fulladder__5_474 genblk1_56_a (.a(x[56]), .b(y[56]), .cin(z[56]), .sum(s1[56]), 
      .carry(c1[56]));
   fulladder__5_482 genblk1_57_a (.a(x[57]), .b(y[57]), .cin(z[57]), .sum(s1[57]), 
      .carry(c1[57]));
   fulladder__5_490 genblk1_58_a (.a(x[63]), .b(y[58]), .cin(z[58]), .sum(s1[58]), 
      .carry(c1[58]));
   fulladder__5_498 genblk1_59_a (.a(x[63]), .b(y[63]), .cin(z[59]), .sum(s1[59]), 
      .carry(c1[59]));
   fulladder__5_506 genblk1_60_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[60]), 
      .carry(c1[60]));
   fulladder__5_514 genblk1_61_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[61]), 
      .carry(c1[61]));
   fulladder__5_522 genblk1_62_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[62]), 
      .carry(c1[62]));
   fulladder__5_530 genblk1_63_a (.a(x[63]), .b(y[63]), .cin(z[63]), .sum(s1[63]), 
      .carry());
   fulladder__5_754 genblk2_28_b (.a(s1[29]), .b(c1[28]), .cin(), .sum(s[29]), 
      .carry(c2[29]));
   fulladder__5_762 genblk2_29_b (.a(s1[30]), .b(c1[29]), .cin(c2[29]), .sum(
      s[30]), .carry(c2[30]));
   fulladder__5_770 genblk2_30_b (.a(s1[31]), .b(c1[30]), .cin(c2[30]), .sum(
      s[31]), .carry(c2[31]));
   fulladder__5_778 genblk2_31_b (.a(s1[32]), .b(c1[31]), .cin(c2[31]), .sum(
      s[32]), .carry(c2[32]));
   fulladder__5_786 genblk2_32_b (.a(s1[33]), .b(c1[32]), .cin(c2[32]), .sum(
      s[33]), .carry(c2[33]));
   fulladder__5_794 genblk2_33_b (.a(s1[34]), .b(c1[33]), .cin(c2[33]), .sum(
      s[34]), .carry(c2[34]));
   fulladder__5_802 genblk2_34_b (.a(s1[35]), .b(c1[34]), .cin(c2[34]), .sum(
      s[35]), .carry(c2[35]));
   fulladder__5_810 genblk2_35_b (.a(s1[36]), .b(c1[35]), .cin(c2[35]), .sum(
      s[36]), .carry(c2[36]));
   fulladder__5_818 genblk2_36_b (.a(s1[37]), .b(c1[36]), .cin(c2[36]), .sum(
      s[37]), .carry(c2[37]));
   fulladder__5_826 genblk2_37_b (.a(s1[38]), .b(c1[37]), .cin(c2[37]), .sum(
      s[38]), .carry(c2[38]));
   fulladder__5_834 genblk2_38_b (.a(s1[39]), .b(c1[38]), .cin(c2[38]), .sum(
      s[39]), .carry(c2[39]));
   fulladder__5_842 genblk2_39_b (.a(s1[40]), .b(c1[39]), .cin(c2[39]), .sum(
      s[40]), .carry(c2[40]));
   fulladder__5_850 genblk2_40_b (.a(s1[41]), .b(c1[40]), .cin(c2[40]), .sum(
      s[41]), .carry(c2[41]));
   fulladder__5_858 genblk2_41_b (.a(s1[42]), .b(c1[41]), .cin(c2[41]), .sum(
      s[42]), .carry(c2[42]));
   fulladder__5_866 genblk2_42_b (.a(s1[43]), .b(c1[42]), .cin(c2[42]), .sum(
      s[43]), .carry(c2[43]));
   fulladder__5_874 genblk2_43_b (.a(s1[44]), .b(c1[43]), .cin(c2[43]), .sum(
      s[44]), .carry(c2[44]));
   fulladder__5_882 genblk2_44_b (.a(s1[45]), .b(c1[44]), .cin(c2[44]), .sum(
      s[45]), .carry(c2[45]));
   fulladder__5_890 genblk2_45_b (.a(s1[46]), .b(c1[45]), .cin(c2[45]), .sum(
      s[46]), .carry(c2[46]));
   fulladder__5_898 genblk2_46_b (.a(s1[47]), .b(c1[46]), .cin(c2[46]), .sum(
      s[47]), .carry(c2[47]));
   fulladder__5_906 genblk2_47_b (.a(s1[48]), .b(c1[47]), .cin(c2[47]), .sum(
      s[48]), .carry(c2[48]));
   fulladder__5_914 genblk2_48_b (.a(s1[49]), .b(c1[48]), .cin(c2[48]), .sum(
      s[49]), .carry(c2[49]));
   fulladder__5_922 genblk2_49_b (.a(s1[50]), .b(c1[49]), .cin(c2[49]), .sum(
      s[50]), .carry(c2[50]));
   fulladder__5_930 genblk2_50_b (.a(s1[51]), .b(c1[50]), .cin(c2[50]), .sum(
      s[51]), .carry(c2[51]));
   fulladder__5_938 genblk2_51_b (.a(s1[52]), .b(c1[51]), .cin(c2[51]), .sum(
      s[52]), .carry(c2[52]));
   fulladder__5_946 genblk2_52_b (.a(s1[53]), .b(c1[52]), .cin(c2[52]), .sum(
      s[53]), .carry(c2[53]));
   fulladder__5_954 genblk2_53_b (.a(s1[54]), .b(c1[53]), .cin(c2[53]), .sum(
      s[54]), .carry(c2[54]));
   fulladder__5_962 genblk2_54_b (.a(s1[55]), .b(c1[54]), .cin(c2[54]), .sum(
      s[55]), .carry(c2[55]));
   fulladder__5_970 genblk2_55_b (.a(s1[56]), .b(c1[55]), .cin(c2[55]), .sum(
      s[56]), .carry(c2[56]));
   fulladder__5_978 genblk2_56_b (.a(s1[57]), .b(c1[56]), .cin(c2[56]), .sum(
      s[57]), .carry(c2[57]));
   fulladder__5_986 genblk2_57_b (.a(s1[58]), .b(c1[57]), .cin(c2[57]), .sum(
      s[58]), .carry(c2[58]));
   fulladder__5_994 genblk2_58_b (.a(s1[59]), .b(c1[58]), .cin(c2[58]), .sum(
      s[59]), .carry(c2[59]));
   fulladder__5_1002 genblk2_59_b (.a(s1[60]), .b(c1[59]), .cin(c2[59]), 
      .sum(s[60]), .carry(c2[60]));
   fulladder__5_1010 genblk2_60_b (.a(s1[61]), .b(c1[60]), .cin(c2[60]), 
      .sum(s[61]), .carry(c2[61]));
   fulladder__5_1018 genblk2_61_b (.a(s1[62]), .b(c1[61]), .cin(c2[61]), 
      .sum(s[62]), .carry(c2[62]));
   fulladder genblk2_62_b (.a(s1[63]), .b(c1[62]), .cin(c2[62]), .sum(s[63]), 
      .carry());
endmodule

module wallace_tree(A, B, Out, clk, rst);
   input [31:0]A;
   input [31:0]B;
   output [63:0]Out;
   input clk;
   input rst;

   wire n_2_10;
   wire n_2_11;
   wire n_2_12;
   wire n_2_13;
   wire n_2_14;
   wire n_2_15;
   wire n_2_16;
   wire n_2_17;
   wire n_2_18;
   wire n_2_19;
   wire n_2_20;
   wire n_2_21;
   wire n_2_22;
   wire n_2_23;
   wire n_2_24;
   wire n_2_25;
   wire n_2_26;
   wire n_2_27;
   wire n_2_28;
   wire n_2_29;
   wire n_2_30;
   wire n_2_31;
   wire n_2_32;
   wire n_2_33;
   wire n_2_34;
   wire n_2_35;
   wire n_2_36;
   wire n_2_37;
   wire n_2_38;
   wire n_2_39;
   wire n_2_40;
   wire n_2_0_0;
   wire n_2_0_1;
   wire n_2_0_2;
   wire n_2_0_3;
   wire n_2_0_4;
   wire n_2_0_5;
   wire n_2_0_6;
   wire n_2_0_7;
   wire n_2_0_8;
   wire n_2_0_9;
   wire n_2_0_10;
   wire n_2_0_11;
   wire n_2_0_12;
   wire n_2_0_13;
   wire n_2_0_14;
   wire n_2_0_15;
   wire n_2_0_16;
   wire n_2_0_17;
   wire n_2_0_18;
   wire n_2_0_19;
   wire n_2_0_20;
   wire n_2_0_21;
   wire n_2_0_22;
   wire n_2_0_23;
   wire n_2_0_24;
   wire n_2_0_25;
   wire n_2_0_26;
   wire n_2_0_27;
   wire n_2_0_28;
   wire n_2_0_29;
   wire n_2_0_30;
   wire n_2_0_31;
   wire n_2_0_32;
   wire n_2_0_33;
   wire n_2_0_34;
   wire n_2_0_35;
   wire n_2_0_36;
   wire n_2_41;
   wire n_2_42;
   wire n_2_43;
   wire n_2_44;
   wire n_2_45;
   wire n_2_46;
   wire n_2_47;
   wire n_2_48;
   wire n_2_49;
   wire n_2_50;
   wire n_2_51;
   wire n_2_52;
   wire n_2_53;
   wire n_2_54;
   wire n_2_55;
   wire n_2_56;
   wire n_2_57;
   wire n_2_58;
   wire n_2_59;
   wire n_2_60;
   wire n_2_61;
   wire n_2_62;
   wire n_2_63;
   wire n_2_64;
   wire n_2_65;
   wire n_2_66;
   wire n_2_67;
   wire n_2_68;
   wire n_2_69;
   wire n_2_70;
   wire n_2_71;
   wire n_2_0_37;
   wire n_2_72;
   wire n_2_73;
   wire n_2_74;
   wire n_2_75;
   wire n_2_76;
   wire n_2_77;
   wire n_2_78;
   wire n_2_79;
   wire n_2_80;
   wire n_2_81;
   wire n_2_82;
   wire n_2_83;
   wire n_2_84;
   wire n_2_85;
   wire n_2_86;
   wire n_2_87;
   wire n_2_88;
   wire n_2_89;
   wire n_2_90;
   wire n_2_91;
   wire n_2_92;
   wire n_2_93;
   wire n_2_94;
   wire n_2_95;
   wire n_2_96;
   wire n_2_97;
   wire n_2_98;
   wire n_2_99;
   wire n_2_100;
   wire n_2_101;
   wire n_2_102;
   wire n_2_103;
   wire n_2_0_38;
   wire n_2_104;
   wire n_2_105;
   wire n_2_106;
   wire n_2_107;
   wire n_2_108;
   wire n_2_109;
   wire n_2_110;
   wire n_2_111;
   wire n_2_112;
   wire n_2_113;
   wire n_2_114;
   wire n_2_115;
   wire n_2_116;
   wire n_2_117;
   wire n_2_118;
   wire n_2_119;
   wire n_2_120;
   wire n_2_121;
   wire n_2_122;
   wire n_2_123;
   wire n_2_124;
   wire n_2_125;
   wire n_2_126;
   wire n_2_127;
   wire n_2_128;
   wire n_2_129;
   wire n_2_130;
   wire n_2_131;
   wire n_2_132;
   wire n_2_133;
   wire n_2_134;
   wire n_2_135;
   wire n_2_0_39;
   wire n_2_136;
   wire n_2_137;
   wire n_2_138;
   wire n_2_139;
   wire n_2_140;
   wire n_2_141;
   wire n_2_142;
   wire n_2_143;
   wire n_2_144;
   wire n_2_145;
   wire n_2_146;
   wire n_2_147;
   wire n_2_148;
   wire n_2_149;
   wire n_2_150;
   wire n_2_151;
   wire n_2_152;
   wire n_2_153;
   wire n_2_154;
   wire n_2_155;
   wire n_2_156;
   wire n_2_157;
   wire n_2_158;
   wire n_2_159;
   wire n_2_160;
   wire n_2_161;
   wire n_2_162;
   wire n_2_163;
   wire n_2_164;
   wire n_2_165;
   wire n_2_166;
   wire n_2_0_40;
   wire n_2_167;
   wire n_2_168;
   wire n_2_169;
   wire n_2_170;
   wire n_2_171;
   wire n_2_172;
   wire n_2_173;
   wire n_2_174;
   wire n_2_175;
   wire n_2_176;
   wire n_2_177;
   wire n_2_178;
   wire n_2_179;
   wire n_2_180;
   wire n_2_181;
   wire n_2_182;
   wire n_2_183;
   wire n_2_184;
   wire n_2_185;
   wire n_2_186;
   wire n_2_187;
   wire n_2_188;
   wire n_2_189;
   wire n_2_190;
   wire n_2_191;
   wire n_2_192;
   wire n_2_193;
   wire n_2_194;
   wire n_2_195;
   wire n_2_196;
   wire n_2_197;
   wire n_2_198;
   wire n_2_0_41;
   wire n_2_199;
   wire n_2_200;
   wire n_2_201;
   wire n_2_202;
   wire n_2_203;
   wire n_2_204;
   wire n_2_205;
   wire n_2_206;
   wire n_2_207;
   wire n_2_208;
   wire n_2_209;
   wire n_2_210;
   wire n_2_211;
   wire n_2_212;
   wire n_2_213;
   wire n_2_214;
   wire n_2_215;
   wire n_2_216;
   wire n_2_217;
   wire n_2_218;
   wire n_2_219;
   wire n_2_220;
   wire n_2_221;
   wire n_2_222;
   wire n_2_223;
   wire n_2_224;
   wire n_2_225;
   wire n_2_226;
   wire n_2_227;
   wire n_2_228;
   wire n_2_229;
   wire n_2_230;
   wire n_2_0_42;
   wire n_2_231;
   wire n_2_232;
   wire n_2_233;
   wire n_2_234;
   wire n_2_235;
   wire n_2_236;
   wire n_2_237;
   wire n_2_238;
   wire n_2_239;
   wire n_2_240;
   wire n_2_241;
   wire n_2_242;
   wire n_2_243;
   wire n_2_244;
   wire n_2_245;
   wire n_2_246;
   wire n_2_247;
   wire n_2_248;
   wire n_2_249;
   wire n_2_250;
   wire n_2_251;
   wire n_2_252;
   wire n_2_253;
   wire n_2_254;
   wire n_2_255;
   wire n_2_256;
   wire n_2_257;
   wire n_2_258;
   wire n_2_259;
   wire n_2_260;
   wire n_2_261;
   wire n_2_0_43;
   wire n_2_262;
   wire n_2_263;
   wire n_2_264;
   wire n_2_265;
   wire n_2_266;
   wire n_2_267;
   wire n_2_268;
   wire n_2_269;
   wire n_2_270;
   wire n_2_271;
   wire n_2_272;
   wire n_2_273;
   wire n_2_274;
   wire n_2_275;
   wire n_2_276;
   wire n_2_277;
   wire n_2_278;
   wire n_2_279;
   wire n_2_280;
   wire n_2_281;
   wire n_2_282;
   wire n_2_283;
   wire n_2_284;
   wire n_2_285;
   wire n_2_286;
   wire n_2_287;
   wire n_2_288;
   wire n_2_289;
   wire n_2_290;
   wire n_2_291;
   wire n_2_292;
   wire n_2_293;
   wire n_2_0_44;
   wire n_2_294;
   wire n_2_295;
   wire n_2_296;
   wire n_2_297;
   wire n_2_298;
   wire n_2_299;
   wire n_2_300;
   wire n_2_301;
   wire n_2_302;
   wire n_2_303;
   wire n_2_304;
   wire n_2_305;
   wire n_2_306;
   wire n_2_307;
   wire n_2_308;
   wire n_2_309;
   wire n_2_310;
   wire n_2_311;
   wire n_2_312;
   wire n_2_313;
   wire n_2_314;
   wire n_2_315;
   wire n_2_316;
   wire n_2_317;
   wire n_2_318;
   wire n_2_319;
   wire n_2_320;
   wire n_2_321;
   wire n_2_322;
   wire n_2_323;
   wire n_2_324;
   wire n_2_325;
   wire n_2_0_45;
   wire n_2_326;
   wire n_2_327;
   wire n_2_328;
   wire n_2_329;
   wire n_2_330;
   wire n_2_331;
   wire n_2_332;
   wire n_2_333;
   wire n_2_334;
   wire n_2_335;
   wire n_2_336;
   wire n_2_337;
   wire n_2_338;
   wire n_2_339;
   wire n_2_340;
   wire n_2_341;
   wire n_2_342;
   wire n_2_343;
   wire n_2_344;
   wire n_2_345;
   wire n_2_346;
   wire n_2_347;
   wire n_2_348;
   wire n_2_349;
   wire n_2_350;
   wire n_2_351;
   wire n_2_352;
   wire n_2_353;
   wire n_2_354;
   wire n_2_355;
   wire n_2_356;
   wire n_2_0_46;
   wire n_2_357;
   wire n_2_358;
   wire n_2_359;
   wire n_2_360;
   wire n_2_361;
   wire n_2_362;
   wire n_2_363;
   wire n_2_364;
   wire n_2_365;
   wire n_2_366;
   wire n_2_367;
   wire n_2_368;
   wire n_2_369;
   wire n_2_370;
   wire n_2_371;
   wire n_2_372;
   wire n_2_373;
   wire n_2_374;
   wire n_2_375;
   wire n_2_376;
   wire n_2_377;
   wire n_2_378;
   wire n_2_379;
   wire n_2_380;
   wire n_2_381;
   wire n_2_382;
   wire n_2_383;
   wire n_2_384;
   wire n_2_385;
   wire n_2_386;
   wire n_2_387;
   wire n_2_388;
   wire n_2_0_47;
   wire n_2_389;
   wire n_2_390;
   wire n_2_391;
   wire n_2_392;
   wire n_2_393;
   wire n_2_394;
   wire n_2_395;
   wire n_2_396;
   wire n_2_397;
   wire n_2_398;
   wire n_2_399;
   wire n_2_400;
   wire n_2_401;
   wire n_2_402;
   wire n_2_403;
   wire n_2_404;
   wire n_2_405;
   wire n_2_406;
   wire n_2_407;
   wire n_2_408;
   wire n_2_409;
   wire n_2_410;
   wire n_2_411;
   wire n_2_412;
   wire n_2_413;
   wire n_2_414;
   wire n_2_415;
   wire n_2_416;
   wire n_2_417;
   wire n_2_418;
   wire n_2_419;
   wire n_2_420;
   wire n_2_0_48;
   wire n_2_421;
   wire n_2_422;
   wire n_2_423;
   wire n_2_424;
   wire n_2_425;
   wire n_2_426;
   wire n_2_427;
   wire n_2_428;
   wire n_2_429;
   wire n_2_430;
   wire n_2_431;
   wire n_2_432;
   wire n_2_433;
   wire n_2_434;
   wire n_2_435;
   wire n_2_436;
   wire n_2_437;
   wire n_2_438;
   wire n_2_439;
   wire n_2_440;
   wire n_2_441;
   wire n_2_442;
   wire n_2_443;
   wire n_2_444;
   wire n_2_445;
   wire n_2_446;
   wire n_2_447;
   wire n_2_448;
   wire n_2_449;
   wire n_2_450;
   wire n_2_451;
   wire n_2_452;
   wire n_2_0_49;
   wire n_2_453;
   wire n_2_454;
   wire n_2_455;
   wire n_2_456;
   wire n_2_457;
   wire n_2_458;
   wire n_2_459;
   wire n_2_460;
   wire n_2_461;
   wire n_2_462;
   wire n_2_463;
   wire n_2_464;
   wire n_2_465;
   wire n_2_466;
   wire n_2_467;
   wire n_2_468;
   wire n_2_469;
   wire n_2_470;
   wire n_2_471;
   wire n_2_472;
   wire n_2_473;
   wire n_2_474;
   wire n_2_475;
   wire n_2_476;
   wire n_2_477;
   wire n_2_478;
   wire n_2_479;
   wire n_2_480;
   wire n_2_481;
   wire n_2_482;
   wire n_2_483;
   wire n_2_484;
   wire n_2_0_50;
   wire n_2_485;
   wire n_2_486;
   wire n_2_487;
   wire n_2_488;
   wire n_2_489;
   wire n_2_490;
   wire n_2_491;
   wire n_2_492;
   wire n_2_493;
   wire n_2_494;
   wire n_2_495;
   wire n_2_496;
   wire n_2_497;
   wire n_2_498;
   wire n_2_499;
   wire n_2_500;
   wire n_2_501;
   wire n_2_502;
   wire n_2_503;
   wire n_2_504;
   wire n_2_505;
   wire n_2_506;
   wire n_2_507;
   wire n_2_508;
   wire n_2_509;
   wire n_2_510;
   wire n_2_511;
   wire n_2_512;
   wire n_2_513;
   wire n_2_514;
   wire n_2_515;
   wire n_2_516;
   wire n_2_0_51;
   wire n_2_517;
   wire n_2_518;
   wire n_2_519;
   wire n_2_520;
   wire n_2_521;
   wire n_2_522;
   wire n_2_523;
   wire n_2_524;
   wire n_2_525;
   wire n_2_526;
   wire n_2_527;
   wire n_2_528;
   wire n_2_529;
   wire n_2_530;
   wire n_2_531;
   wire n_2_532;
   wire n_2_533;
   wire n_2_534;
   wire n_2_535;
   wire n_2_536;
   wire n_2_537;
   wire n_2_538;
   wire n_2_539;
   wire n_2_540;
   wire n_2_541;
   wire n_2_542;
   wire n_2_543;
   wire n_2_544;
   wire n_2_545;
   wire n_2_546;
   wire n_2_547;
   wire n_2_548;
   wire n_2_0_52;
   wire n_2_549;
   wire n_2_550;
   wire n_2_551;
   wire n_2_552;
   wire n_2_553;
   wire n_2_554;
   wire n_2_555;
   wire n_2_556;
   wire n_2_557;
   wire n_2_558;
   wire n_2_559;
   wire n_2_560;
   wire n_2_561;
   wire n_2_562;
   wire n_2_563;
   wire n_2_564;
   wire n_2_565;
   wire n_2_566;
   wire n_2_567;
   wire n_2_568;
   wire n_2_569;
   wire n_2_570;
   wire n_2_571;
   wire n_2_572;
   wire n_2_573;
   wire n_2_574;
   wire n_2_575;
   wire n_2_576;
   wire n_2_577;
   wire n_2_578;
   wire n_2_579;
   wire n_2_580;
   wire n_2_0_53;
   wire n_2_581;
   wire n_2_582;
   wire n_2_583;
   wire n_2_584;
   wire n_2_585;
   wire n_2_586;
   wire n_2_587;
   wire n_2_588;
   wire n_2_589;
   wire n_2_590;
   wire n_2_591;
   wire n_2_592;
   wire n_2_593;
   wire n_2_594;
   wire n_2_595;
   wire n_2_596;
   wire n_2_597;
   wire n_2_598;
   wire n_2_599;
   wire n_2_600;
   wire n_2_601;
   wire n_2_602;
   wire n_2_603;
   wire n_2_604;
   wire n_2_605;
   wire n_2_606;
   wire n_2_607;
   wire n_2_608;
   wire n_2_609;
   wire n_2_610;
   wire n_2_611;
   wire n_2_612;
   wire n_2_0_54;
   wire n_2_613;
   wire n_2_614;
   wire n_2_615;
   wire n_2_616;
   wire n_2_617;
   wire n_2_618;
   wire n_2_619;
   wire n_2_620;
   wire n_2_621;
   wire n_2_622;
   wire n_2_623;
   wire n_2_624;
   wire n_2_625;
   wire n_2_626;
   wire n_2_627;
   wire n_2_628;
   wire n_2_629;
   wire n_2_630;
   wire n_2_631;
   wire n_2_632;
   wire n_2_633;
   wire n_2_634;
   wire n_2_635;
   wire n_2_636;
   wire n_2_637;
   wire n_2_638;
   wire n_2_639;
   wire n_2_640;
   wire n_2_641;
   wire n_2_642;
   wire n_2_643;
   wire n_2_0_55;
   wire n_2_644;
   wire n_2_645;
   wire n_2_646;
   wire n_2_647;
   wire n_2_648;
   wire n_2_649;
   wire n_2_650;
   wire n_2_651;
   wire n_2_652;
   wire n_2_653;
   wire n_2_654;
   wire n_2_655;
   wire n_2_656;
   wire n_2_657;
   wire n_2_658;
   wire n_2_659;
   wire n_2_660;
   wire n_2_661;
   wire n_2_662;
   wire n_2_663;
   wire n_2_664;
   wire n_2_665;
   wire n_2_666;
   wire n_2_667;
   wire n_2_668;
   wire n_2_669;
   wire n_2_670;
   wire n_2_671;
   wire n_2_672;
   wire n_2_673;
   wire n_2_674;
   wire n_2_675;
   wire n_2_0_56;
   wire n_2_676;
   wire n_2_677;
   wire n_2_678;
   wire n_2_679;
   wire n_2_680;
   wire n_2_681;
   wire n_2_682;
   wire n_2_683;
   wire n_2_684;
   wire n_2_685;
   wire n_2_686;
   wire n_2_687;
   wire n_2_688;
   wire n_2_689;
   wire n_2_690;
   wire n_2_691;
   wire n_2_692;
   wire n_2_693;
   wire n_2_694;
   wire n_2_695;
   wire n_2_696;
   wire n_2_697;
   wire n_2_698;
   wire n_2_699;
   wire n_2_700;
   wire n_2_701;
   wire n_2_702;
   wire n_2_712;
   wire n_2_713__0;
   wire n_2_714__0;
   wire n_2_779;
   wire n_2_846;
   wire n_2_0_57;
   wire n_2_0_58;
   wire n_2_0_59;
   wire n_2_0_60;
   wire n_2_0_61;
   wire n_2_0_62;
   wire n_2_713__1;
   wire n_2_714__1;
   wire n_2_715;
   wire n_2_716;
   wire n_2_717;
   wire n_2_718;
   wire n_2_719;
   wire n_2_720;
   wire n_2_721;
   wire n_2_722;
   wire n_2_723;
   wire n_2_724;
   wire n_2_725;
   wire n_2_726;
   wire n_2_727;
   wire n_2_728;
   wire n_2_729;
   wire n_2_730;
   wire n_2_731;
   wire n_2_732;
   wire n_2_733;
   wire n_2_734;
   wire n_2_735;
   wire n_2_736;
   wire n_2_737;
   wire n_2_738;
   wire n_2_739;
   wire n_2_740;
   wire n_2_741;
   wire n_2_742;
   wire n_2_743;
   wire n_2_744;
   wire n_2_745;
   wire n_2_746;
   wire n_2_747;
   wire n_2_748;
   wire n_2_749;
   wire n_2_750;
   wire n_2_751;
   wire n_2_752;
   wire n_2_753;
   wire n_2_754;
   wire n_2_755;
   wire n_2_756;
   wire n_2_757;
   wire n_2_758;
   wire n_2_759;
   wire n_2_760;
   wire n_2_761;
   wire n_2_762;
   wire n_2_763;
   wire n_2_764;
   wire n_2_765;
   wire n_2_766;
   wire n_2_780;
   wire n_2_781;
   wire n_2_782;
   wire n_2_783;
   wire n_2_784;
   wire n_2_785;
   wire n_2_786;
   wire n_2_787;
   wire n_2_788;
   wire n_2_789;
   wire n_2_790;
   wire n_2_791;
   wire n_2_792;
   wire n_2_793;
   wire n_2_794;
   wire n_2_795;
   wire n_2_796;
   wire n_2_797;
   wire n_2_798;
   wire n_2_799;
   wire n_2_800;
   wire n_2_801;
   wire n_2_802;
   wire n_2_803;
   wire n_2_804;
   wire n_2_805;
   wire n_2_806;
   wire n_2_807;
   wire n_2_808;
   wire n_2_809;
   wire n_2_810;
   wire n_2_811;
   wire n_2_812;
   wire n_2_813;
   wire n_2_814;
   wire n_2_815;
   wire n_2_816;
   wire n_2_817;
   wire n_2_818;
   wire n_2_819;
   wire n_2_820;
   wire n_2_821;
   wire n_2_822;
   wire n_2_823;
   wire n_2_824;
   wire n_2_825;
   wire n_2_826;
   wire n_2_827;
   wire n_2_828;
   wire n_2_829;
   wire n_2_830;
   wire n_2_847;
   wire n_2_848;
   wire n_2_0;
   wire n_2_1;
   wire n_2_2;
   wire n_2_3;
   wire n_2_4;
   wire n_2_5;
   wire n_2_6;
   wire n_2_7;
   wire n_2_8;
   wire n_2_9;
   wire n_2_703;
   wire n_2_704;
   wire n_2_705;
   wire n_2_706;
   wire n_2_707;
   wire n_2_708;
   wire n_2_709;
   wire n_2_710;
   wire n_2_711;
   wire n_2_767;
   wire n_2_768;
   wire n_2_769;
   wire n_2_770;
   wire n_2_771;
   wire n_2_772;
   wire n_2_773;
   wire n_2_774;
   wire n_2_775;
   wire n_2_776;
   wire n_2_777;
   wire n_2_778;
   wire n_2_831;
   wire n_2_832;
   wire n_2_833;
   wire n_2_834;
   wire n_2_835;
   wire n_2_836;
   wire n_2_837;
   wire n_2_838;
   wire n_2_839;
   wire n_2_840;
   wire n_2_841;
   wire n_2_842;
   wire n_2_843;
   wire n_2_844;
   wire n_2_845;
   wire n_5_22;
   wire n_5_23;
   wire n_5_24;
   wire n_5_25;
   wire n_5_26;
   wire n_5_27;
   wire n_5_28;
   wire n_5_29;
   wire n_5_30;
   wire n_5_31;
   wire n_5_32;
   wire n_5_33;
   wire n_5_34;
   wire n_5_35;
   wire n_5_36;
   wire n_5_37;
   wire n_5_38;
   wire n_5_39;
   wire n_5_40;
   wire n_5_41;
   wire n_5_42;
   wire n_5_43;
   wire n_5_44;
   wire n_5_45;
   wire n_5_46;
   wire n_5_47;
   wire n_5_48;
   wire n_5_49;
   wire n_5_50;
   wire n_5_51;
   wire n_5_52;
   wire n_5_53;
   wire n_5_54;
   wire n_5_55;
   wire n_5_56;
   wire n_5_57;
   wire n_5_58;
   wire n_5_59;
   wire n_5_60;
   wire n_5_61;
   wire n_5_62;
   wire n_5_63;
   wire n_5_0;
   wire n_5_1;
   wire n_5_2;
   wire n_5_3;
   wire n_5_4;
   wire n_5_5;
   wire n_5_6;
   wire n_5_7;
   wire n_5_8;
   wire n_5_9;
   wire n_5_10;
   wire n_5_11;
   wire n_5_12;
   wire n_5_13;
   wire n_5_14;
   wire n_5_15;
   wire n_5_16;
   wire n_5_17;
   wire n_5_18;
   wire n_5_19;
   wire n_5_20;
   wire n_5_21;
   wire n_5_64;
   wire n_5_65;
   wire n_5_66;
   wire n_5_67;
   wire n_5_68;
   wire n_5_69;
   wire n_5_70;
   wire n_5_71;
   wire n_5_72;
   wire n_5_73;
   wire n_5_74;
   wire n_5_75;
   wire n_5_76;
   wire n_5_77;
   wire n_5_78;
   wire n_5_79;
   wire n_5_80;
   wire n_5_81;
   wire n_5_82;
   wire n_5_83;
   wire n_5_84;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire [63:0]product;
   wire y;
   wire [31:0]x;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_128;
   wire n_0_129;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_64;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;

   datapath i_2_27 (.p_0({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, 
      uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, 
      uc_30, uc_31, n_2_40, n_2_39, n_2_38, n_2_37, n_2_36, n_2_35, n_2_34, 
      n_2_33, n_2_32, n_2_31, n_2_30, n_2_29, n_2_28, n_2_27, n_2_26, n_2_25, 
      n_2_24, n_2_23, n_2_22, n_2_21, n_2_20, n_2_19, n_2_18, n_2_17, n_2_16, 
      n_2_15, n_2_14, n_2_13, n_2_12, n_2_11, n_2_10, uc_32}), .p_1({1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, x[31], x[30], x[29], x[28], x[27], 
      x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], 
      x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], 
      x[5], x[4], x[3], x[2], x[1], x[0]}));
   INV_X1 i_2_0_0 (.A(n_819), .ZN(n_2_0_0));
   INV_X1 i_2_0_1 (.A(x[0]), .ZN(n_2_0_1));
   NOR2_X1 i_2_0_2 (.A1(n_2_0_0), .A2(n_2_0_1), .ZN(n_0));
   INV_X1 i_2_0_3 (.A(x[1]), .ZN(n_2_0_2));
   NOR2_X1 i_2_0_4 (.A1(n_2_0_0), .A2(n_2_0_2), .ZN(n_1));
   INV_X1 i_2_0_5 (.A(x[2]), .ZN(n_2_0_3));
   NOR2_X1 i_2_0_6 (.A1(n_2_0_0), .A2(n_2_0_3), .ZN(n_2));
   INV_X1 i_2_0_7 (.A(x[3]), .ZN(n_2_0_4));
   NOR2_X1 i_2_0_8 (.A1(n_2_0_0), .A2(n_2_0_4), .ZN(n_3));
   INV_X1 i_2_0_9 (.A(x[4]), .ZN(n_2_0_5));
   NOR2_X1 i_2_0_10 (.A1(n_2_0_0), .A2(n_2_0_5), .ZN(n_4));
   INV_X1 i_2_0_11 (.A(x[5]), .ZN(n_2_0_6));
   NOR2_X1 i_2_0_12 (.A1(n_2_0_0), .A2(n_2_0_6), .ZN(n_5));
   INV_X1 i_2_0_13 (.A(x[6]), .ZN(n_2_0_7));
   NOR2_X1 i_2_0_14 (.A1(n_2_0_0), .A2(n_2_0_7), .ZN(n_6));
   INV_X1 i_2_0_15 (.A(x[7]), .ZN(n_2_0_8));
   NOR2_X1 i_2_0_16 (.A1(n_2_0_0), .A2(n_2_0_8), .ZN(n_7));
   INV_X1 i_2_0_17 (.A(x[8]), .ZN(n_2_0_9));
   NOR2_X1 i_2_0_18 (.A1(n_2_0_0), .A2(n_2_0_9), .ZN(n_8));
   INV_X1 i_2_0_19 (.A(x[9]), .ZN(n_2_0_10));
   NOR2_X1 i_2_0_20 (.A1(n_2_0_0), .A2(n_2_0_10), .ZN(n_9));
   INV_X1 i_2_0_21 (.A(x[10]), .ZN(n_2_0_11));
   NOR2_X1 i_2_0_22 (.A1(n_2_0_0), .A2(n_2_0_11), .ZN(n_10));
   INV_X1 i_2_0_23 (.A(x[11]), .ZN(n_2_0_12));
   NOR2_X1 i_2_0_24 (.A1(n_2_0_0), .A2(n_2_0_12), .ZN(n_11));
   INV_X1 i_2_0_25 (.A(x[12]), .ZN(n_2_0_13));
   NOR2_X1 i_2_0_26 (.A1(n_2_0_0), .A2(n_2_0_13), .ZN(n_12));
   INV_X1 i_2_0_27 (.A(x[13]), .ZN(n_2_0_14));
   NOR2_X1 i_2_0_28 (.A1(n_2_0_0), .A2(n_2_0_14), .ZN(n_13));
   INV_X1 i_2_0_29 (.A(x[14]), .ZN(n_2_0_15));
   NOR2_X1 i_2_0_30 (.A1(n_2_0_0), .A2(n_2_0_15), .ZN(n_14));
   INV_X1 i_2_0_31 (.A(x[15]), .ZN(n_2_0_16));
   NOR2_X1 i_2_0_32 (.A1(n_2_0_0), .A2(n_2_0_16), .ZN(n_15));
   INV_X1 i_2_0_33 (.A(x[16]), .ZN(n_2_0_17));
   NOR2_X1 i_2_0_34 (.A1(n_2_0_0), .A2(n_2_0_17), .ZN(n_16));
   INV_X1 i_2_0_35 (.A(x[17]), .ZN(n_2_0_18));
   NOR2_X1 i_2_0_36 (.A1(n_2_0_0), .A2(n_2_0_18), .ZN(n_17));
   INV_X1 i_2_0_37 (.A(x[18]), .ZN(n_2_0_19));
   NOR2_X1 i_2_0_38 (.A1(n_2_0_0), .A2(n_2_0_19), .ZN(n_18));
   INV_X1 i_2_0_39 (.A(x[19]), .ZN(n_2_0_20));
   NOR2_X1 i_2_0_40 (.A1(n_2_0_0), .A2(n_2_0_20), .ZN(n_19));
   INV_X1 i_2_0_41 (.A(x[20]), .ZN(n_2_0_21));
   NOR2_X1 i_2_0_42 (.A1(n_2_0_0), .A2(n_2_0_21), .ZN(n_20));
   INV_X1 i_2_0_43 (.A(x[21]), .ZN(n_2_0_22));
   NOR2_X1 i_2_0_44 (.A1(n_2_0_0), .A2(n_2_0_22), .ZN(n_21));
   INV_X1 i_2_0_45 (.A(x[22]), .ZN(n_2_0_23));
   NOR2_X1 i_2_0_46 (.A1(n_2_0_0), .A2(n_2_0_23), .ZN(n_22));
   INV_X1 i_2_0_47 (.A(x[23]), .ZN(n_2_0_24));
   NOR2_X1 i_2_0_48 (.A1(n_2_0_0), .A2(n_2_0_24), .ZN(n_23));
   INV_X1 i_2_0_49 (.A(x[24]), .ZN(n_2_0_25));
   NOR2_X1 i_2_0_50 (.A1(n_2_0_0), .A2(n_2_0_25), .ZN(n_24));
   INV_X1 i_2_0_51 (.A(x[25]), .ZN(n_2_0_26));
   NOR2_X1 i_2_0_52 (.A1(n_2_0_0), .A2(n_2_0_26), .ZN(n_25));
   INV_X1 i_2_0_53 (.A(x[26]), .ZN(n_2_0_27));
   NOR2_X1 i_2_0_54 (.A1(n_2_0_0), .A2(n_2_0_27), .ZN(n_26));
   INV_X1 i_2_0_55 (.A(x[27]), .ZN(n_2_0_28));
   NOR2_X1 i_2_0_56 (.A1(n_2_0_0), .A2(n_2_0_28), .ZN(n_27));
   INV_X1 i_2_0_57 (.A(x[28]), .ZN(n_2_0_29));
   NOR2_X1 i_2_0_58 (.A1(n_2_0_0), .A2(n_2_0_29), .ZN(n_28));
   INV_X1 i_2_0_59 (.A(x[29]), .ZN(n_2_0_30));
   NOR2_X1 i_2_0_60 (.A1(n_2_0_0), .A2(n_2_0_30), .ZN(n_29));
   INV_X1 i_2_0_61 (.A(x[30]), .ZN(n_2_0_31));
   NOR2_X1 i_2_0_62 (.A1(n_2_0_0), .A2(n_2_0_31), .ZN(n_30));
   INV_X1 i_2_0_63 (.A(x[31]), .ZN(n_2_0_32));
   NOR2_X1 i_2_0_64 (.A1(n_2_0_0), .A2(n_2_0_32), .ZN(n_31));
   INV_X1 i_2_0_65 (.A(n_818), .ZN(n_2_0_33));
   NOR2_X1 i_2_0_66 (.A1(n_2_0_33), .A2(n_2_0_1), .ZN(n_32));
   NOR2_X1 i_2_0_67 (.A1(n_2_0_33), .A2(n_2_0_2), .ZN(n_33));
   NOR2_X1 i_2_0_68 (.A1(n_2_0_33), .A2(n_2_0_3), .ZN(n_34));
   NOR2_X1 i_2_0_69 (.A1(n_2_0_33), .A2(n_2_0_4), .ZN(n_35));
   NOR2_X1 i_2_0_70 (.A1(n_2_0_33), .A2(n_2_0_5), .ZN(n_36));
   NOR2_X1 i_2_0_71 (.A1(n_2_0_33), .A2(n_2_0_6), .ZN(n_37));
   NOR2_X1 i_2_0_72 (.A1(n_2_0_33), .A2(n_2_0_7), .ZN(n_38));
   NOR2_X1 i_2_0_73 (.A1(n_2_0_33), .A2(n_2_0_8), .ZN(n_39));
   NOR2_X1 i_2_0_74 (.A1(n_2_0_33), .A2(n_2_0_9), .ZN(n_40));
   NOR2_X1 i_2_0_75 (.A1(n_2_0_33), .A2(n_2_0_10), .ZN(n_41));
   NOR2_X1 i_2_0_76 (.A1(n_2_0_33), .A2(n_2_0_11), .ZN(n_42));
   NOR2_X1 i_2_0_77 (.A1(n_2_0_33), .A2(n_2_0_12), .ZN(n_43));
   NOR2_X1 i_2_0_78 (.A1(n_2_0_33), .A2(n_2_0_13), .ZN(n_44));
   NOR2_X1 i_2_0_79 (.A1(n_2_0_33), .A2(n_2_0_14), .ZN(n_45));
   NOR2_X1 i_2_0_80 (.A1(n_2_0_33), .A2(n_2_0_15), .ZN(n_46));
   NOR2_X1 i_2_0_81 (.A1(n_2_0_33), .A2(n_2_0_16), .ZN(n_47));
   NOR2_X1 i_2_0_82 (.A1(n_2_0_33), .A2(n_2_0_17), .ZN(n_48));
   NOR2_X1 i_2_0_83 (.A1(n_2_0_33), .A2(n_2_0_18), .ZN(n_49));
   NOR2_X1 i_2_0_84 (.A1(n_2_0_33), .A2(n_2_0_19), .ZN(n_50));
   NOR2_X1 i_2_0_85 (.A1(n_2_0_33), .A2(n_2_0_20), .ZN(n_51));
   NOR2_X1 i_2_0_86 (.A1(n_2_0_33), .A2(n_2_0_21), .ZN(n_52));
   NOR2_X1 i_2_0_87 (.A1(n_2_0_33), .A2(n_2_0_22), .ZN(n_53));
   NOR2_X1 i_2_0_88 (.A1(n_2_0_33), .A2(n_2_0_23), .ZN(n_54));
   NOR2_X1 i_2_0_89 (.A1(n_2_0_33), .A2(n_2_0_24), .ZN(n_55));
   NOR2_X1 i_2_0_90 (.A1(n_2_0_33), .A2(n_2_0_25), .ZN(n_56));
   NOR2_X1 i_2_0_91 (.A1(n_2_0_33), .A2(n_2_0_26), .ZN(n_57));
   NOR2_X1 i_2_0_92 (.A1(n_2_0_33), .A2(n_2_0_27), .ZN(n_58));
   NOR2_X1 i_2_0_93 (.A1(n_2_0_33), .A2(n_2_0_28), .ZN(n_59));
   NOR2_X1 i_2_0_94 (.A1(n_2_0_33), .A2(n_2_0_29), .ZN(n_60));
   NOR2_X1 i_2_0_95 (.A1(n_2_0_33), .A2(n_2_0_30), .ZN(n_61));
   NOR2_X1 i_2_0_96 (.A1(n_2_0_33), .A2(n_2_0_31), .ZN(n_62));
   NOR2_X1 i_2_0_97 (.A1(n_2_0_33), .A2(n_2_0_32), .ZN(n_63));
   INV_X1 i_2_0_98 (.A(n_817), .ZN(n_2_0_34));
   NOR2_X1 i_2_0_99 (.A1(n_2_0_34), .A2(n_2_0_1), .ZN(n_64));
   NOR2_X1 i_2_0_100 (.A1(n_2_0_34), .A2(n_2_0_2), .ZN(n_65));
   NOR2_X1 i_2_0_101 (.A1(n_2_0_34), .A2(n_2_0_3), .ZN(n_66));
   NOR2_X1 i_2_0_102 (.A1(n_2_0_34), .A2(n_2_0_4), .ZN(n_67));
   NOR2_X1 i_2_0_103 (.A1(n_2_0_34), .A2(n_2_0_5), .ZN(n_68));
   NOR2_X1 i_2_0_104 (.A1(n_2_0_34), .A2(n_2_0_6), .ZN(n_69));
   NOR2_X1 i_2_0_105 (.A1(n_2_0_34), .A2(n_2_0_7), .ZN(n_70));
   NOR2_X1 i_2_0_106 (.A1(n_2_0_34), .A2(n_2_0_8), .ZN(n_71));
   NOR2_X1 i_2_0_107 (.A1(n_2_0_34), .A2(n_2_0_9), .ZN(n_72));
   NOR2_X1 i_2_0_108 (.A1(n_2_0_34), .A2(n_2_0_10), .ZN(n_73));
   NOR2_X1 i_2_0_109 (.A1(n_2_0_34), .A2(n_2_0_11), .ZN(n_74));
   NOR2_X1 i_2_0_110 (.A1(n_2_0_34), .A2(n_2_0_12), .ZN(n_75));
   NOR2_X1 i_2_0_111 (.A1(n_2_0_34), .A2(n_2_0_13), .ZN(n_76));
   NOR2_X1 i_2_0_112 (.A1(n_2_0_34), .A2(n_2_0_14), .ZN(n_77));
   NOR2_X1 i_2_0_113 (.A1(n_2_0_34), .A2(n_2_0_15), .ZN(n_78));
   NOR2_X1 i_2_0_114 (.A1(n_2_0_34), .A2(n_2_0_16), .ZN(n_79));
   NOR2_X1 i_2_0_115 (.A1(n_2_0_34), .A2(n_2_0_17), .ZN(n_80));
   NOR2_X1 i_2_0_116 (.A1(n_2_0_34), .A2(n_2_0_18), .ZN(n_81));
   NOR2_X1 i_2_0_117 (.A1(n_2_0_34), .A2(n_2_0_19), .ZN(n_82));
   NOR2_X1 i_2_0_118 (.A1(n_2_0_34), .A2(n_2_0_20), .ZN(n_83));
   NOR2_X1 i_2_0_119 (.A1(n_2_0_34), .A2(n_2_0_21), .ZN(n_84));
   NOR2_X1 i_2_0_120 (.A1(n_2_0_34), .A2(n_2_0_22), .ZN(n_85));
   NOR2_X1 i_2_0_121 (.A1(n_2_0_34), .A2(n_2_0_23), .ZN(n_86));
   NOR2_X1 i_2_0_122 (.A1(n_2_0_34), .A2(n_2_0_24), .ZN(n_87));
   NOR2_X1 i_2_0_123 (.A1(n_2_0_34), .A2(n_2_0_25), .ZN(n_88));
   NOR2_X1 i_2_0_124 (.A1(n_2_0_34), .A2(n_2_0_26), .ZN(n_89));
   NOR2_X1 i_2_0_125 (.A1(n_2_0_34), .A2(n_2_0_27), .ZN(n_90));
   NOR2_X1 i_2_0_126 (.A1(n_2_0_34), .A2(n_2_0_28), .ZN(n_91));
   NOR2_X1 i_2_0_127 (.A1(n_2_0_34), .A2(n_2_0_29), .ZN(n_92));
   NOR2_X1 i_2_0_128 (.A1(n_2_0_34), .A2(n_2_0_30), .ZN(n_93));
   NOR2_X1 i_2_0_129 (.A1(n_2_0_34), .A2(n_2_0_31), .ZN(n_94));
   NOR2_X1 i_2_0_130 (.A1(n_2_0_34), .A2(n_2_0_32), .ZN(n_95));
   INV_X1 i_2_0_131 (.A(n_816), .ZN(n_2_0_35));
   NOR2_X1 i_2_0_132 (.A1(n_2_0_35), .A2(n_2_0_1), .ZN(n_96));
   NOR2_X1 i_2_0_133 (.A1(n_2_0_35), .A2(n_2_0_2), .ZN(n_97));
   NOR2_X1 i_2_0_134 (.A1(n_2_0_35), .A2(n_2_0_3), .ZN(n_98));
   NOR2_X1 i_2_0_135 (.A1(n_2_0_35), .A2(n_2_0_4), .ZN(n_99));
   NOR2_X1 i_2_0_136 (.A1(n_2_0_35), .A2(n_2_0_5), .ZN(n_100));
   NOR2_X1 i_2_0_137 (.A1(n_2_0_35), .A2(n_2_0_6), .ZN(n_101));
   NOR2_X1 i_2_0_138 (.A1(n_2_0_35), .A2(n_2_0_7), .ZN(n_102));
   NOR2_X1 i_2_0_139 (.A1(n_2_0_35), .A2(n_2_0_8), .ZN(n_103));
   NOR2_X1 i_2_0_140 (.A1(n_2_0_35), .A2(n_2_0_9), .ZN(n_104));
   NOR2_X1 i_2_0_141 (.A1(n_2_0_35), .A2(n_2_0_10), .ZN(n_105));
   NOR2_X1 i_2_0_142 (.A1(n_2_0_35), .A2(n_2_0_11), .ZN(n_106));
   NOR2_X1 i_2_0_143 (.A1(n_2_0_35), .A2(n_2_0_12), .ZN(n_107));
   NOR2_X1 i_2_0_144 (.A1(n_2_0_35), .A2(n_2_0_13), .ZN(n_108));
   NOR2_X1 i_2_0_145 (.A1(n_2_0_35), .A2(n_2_0_14), .ZN(n_109));
   NOR2_X1 i_2_0_146 (.A1(n_2_0_35), .A2(n_2_0_15), .ZN(n_110));
   NOR2_X1 i_2_0_147 (.A1(n_2_0_35), .A2(n_2_0_16), .ZN(n_111));
   NOR2_X1 i_2_0_148 (.A1(n_2_0_35), .A2(n_2_0_17), .ZN(n_112));
   NOR2_X1 i_2_0_149 (.A1(n_2_0_35), .A2(n_2_0_18), .ZN(n_113));
   NOR2_X1 i_2_0_150 (.A1(n_2_0_35), .A2(n_2_0_19), .ZN(n_114));
   NOR2_X1 i_2_0_151 (.A1(n_2_0_35), .A2(n_2_0_20), .ZN(n_115));
   NOR2_X1 i_2_0_152 (.A1(n_2_0_35), .A2(n_2_0_21), .ZN(n_116));
   NOR2_X1 i_2_0_153 (.A1(n_2_0_35), .A2(n_2_0_22), .ZN(n_117));
   NOR2_X1 i_2_0_154 (.A1(n_2_0_35), .A2(n_2_0_23), .ZN(n_118));
   NOR2_X1 i_2_0_155 (.A1(n_2_0_35), .A2(n_2_0_24), .ZN(n_119));
   NOR2_X1 i_2_0_156 (.A1(n_2_0_35), .A2(n_2_0_25), .ZN(n_120));
   NOR2_X1 i_2_0_157 (.A1(n_2_0_35), .A2(n_2_0_26), .ZN(n_121));
   NOR2_X1 i_2_0_158 (.A1(n_2_0_35), .A2(n_2_0_27), .ZN(n_122));
   NOR2_X1 i_2_0_159 (.A1(n_2_0_35), .A2(n_2_0_28), .ZN(n_123));
   NOR2_X1 i_2_0_160 (.A1(n_2_0_35), .A2(n_2_0_29), .ZN(n_124));
   NOR2_X1 i_2_0_161 (.A1(n_2_0_35), .A2(n_2_0_30), .ZN(n_125));
   NOR2_X1 i_2_0_162 (.A1(n_2_0_35), .A2(n_2_0_31), .ZN(n_126));
   NOR2_X1 i_2_0_163 (.A1(n_2_0_35), .A2(n_2_0_32), .ZN(n_127));
   AND2_X1 i_2_0_164 (.A1(n_815), .A2(x[0]), .ZN(n_128));
   AND2_X1 i_2_0_165 (.A1(n_2_10), .A2(n_815), .ZN(n_129));
   AND2_X1 i_2_0_166 (.A1(n_2_11), .A2(n_815), .ZN(n_130));
   AND2_X1 i_2_0_167 (.A1(n_2_12), .A2(n_815), .ZN(n_131));
   AND2_X1 i_2_0_168 (.A1(n_2_13), .A2(n_815), .ZN(n_132));
   AND2_X1 i_2_0_169 (.A1(n_2_14), .A2(n_815), .ZN(n_133));
   AND2_X1 i_2_0_170 (.A1(n_2_15), .A2(n_815), .ZN(n_134));
   AND2_X1 i_2_0_171 (.A1(n_2_16), .A2(n_815), .ZN(n_135));
   AND2_X1 i_2_0_172 (.A1(n_2_17), .A2(n_815), .ZN(n_136));
   AND2_X1 i_2_0_173 (.A1(n_2_18), .A2(n_815), .ZN(n_137));
   AND2_X1 i_2_0_174 (.A1(n_2_19), .A2(n_815), .ZN(n_138));
   AND2_X1 i_2_0_175 (.A1(n_2_20), .A2(n_815), .ZN(n_139));
   AND2_X1 i_2_0_176 (.A1(n_2_21), .A2(n_815), .ZN(n_140));
   AND2_X1 i_2_0_177 (.A1(n_2_22), .A2(n_815), .ZN(n_141));
   AND2_X1 i_2_0_178 (.A1(n_2_23), .A2(n_815), .ZN(n_142));
   AND2_X1 i_2_0_179 (.A1(n_2_24), .A2(n_815), .ZN(n_143));
   AND2_X1 i_2_0_180 (.A1(n_2_25), .A2(n_815), .ZN(n_144));
   AND2_X1 i_2_0_181 (.A1(n_2_26), .A2(n_815), .ZN(n_145));
   AND2_X1 i_2_0_182 (.A1(n_2_27), .A2(n_815), .ZN(n_146));
   AND2_X1 i_2_0_183 (.A1(n_2_28), .A2(n_815), .ZN(n_147));
   AND2_X1 i_2_0_184 (.A1(n_2_29), .A2(n_815), .ZN(n_148));
   AND2_X1 i_2_0_185 (.A1(n_2_30), .A2(n_815), .ZN(n_149));
   AND2_X1 i_2_0_186 (.A1(n_2_31), .A2(n_815), .ZN(n_150));
   AND2_X1 i_2_0_187 (.A1(n_2_32), .A2(n_815), .ZN(n_151));
   AND2_X1 i_2_0_188 (.A1(n_2_33), .A2(n_815), .ZN(n_152));
   AND2_X1 i_2_0_189 (.A1(n_2_34), .A2(n_815), .ZN(n_153));
   AND2_X1 i_2_0_190 (.A1(n_2_35), .A2(n_815), .ZN(n_154));
   AND2_X1 i_2_0_191 (.A1(n_2_36), .A2(n_815), .ZN(n_155));
   AND2_X1 i_2_0_192 (.A1(n_2_37), .A2(n_815), .ZN(n_156));
   AND2_X1 i_2_0_193 (.A1(n_2_38), .A2(n_815), .ZN(n_157));
   AND2_X1 i_2_0_194 (.A1(n_2_39), .A2(n_815), .ZN(n_158));
   AND2_X1 i_2_0_195 (.A1(n_2_40), .A2(n_815), .ZN(n_159));
   INV_X1 i_2_0_196 (.A(n_814), .ZN(n_2_0_36));
   NOR2_X1 i_2_0_197 (.A1(n_2_0_36), .A2(n_2_0_1), .ZN(n_160));
   NOR2_X1 i_2_0_198 (.A1(n_2_0_36), .A2(n_2_0_2), .ZN(n_2_41));
   NOR2_X1 i_2_0_199 (.A1(n_2_0_36), .A2(n_2_0_3), .ZN(n_2_42));
   NOR2_X1 i_2_0_200 (.A1(n_2_0_36), .A2(n_2_0_4), .ZN(n_2_43));
   NOR2_X1 i_2_0_201 (.A1(n_2_0_36), .A2(n_2_0_5), .ZN(n_2_44));
   NOR2_X1 i_2_0_202 (.A1(n_2_0_36), .A2(n_2_0_6), .ZN(n_2_45));
   NOR2_X1 i_2_0_203 (.A1(n_2_0_36), .A2(n_2_0_7), .ZN(n_2_46));
   NOR2_X1 i_2_0_204 (.A1(n_2_0_36), .A2(n_2_0_8), .ZN(n_2_47));
   NOR2_X1 i_2_0_205 (.A1(n_2_0_36), .A2(n_2_0_9), .ZN(n_2_48));
   NOR2_X1 i_2_0_206 (.A1(n_2_0_36), .A2(n_2_0_10), .ZN(n_2_49));
   NOR2_X1 i_2_0_207 (.A1(n_2_0_36), .A2(n_2_0_11), .ZN(n_2_50));
   NOR2_X1 i_2_0_208 (.A1(n_2_0_36), .A2(n_2_0_12), .ZN(n_2_51));
   NOR2_X1 i_2_0_209 (.A1(n_2_0_36), .A2(n_2_0_13), .ZN(n_2_52));
   NOR2_X1 i_2_0_210 (.A1(n_2_0_36), .A2(n_2_0_14), .ZN(n_2_53));
   NOR2_X1 i_2_0_211 (.A1(n_2_0_36), .A2(n_2_0_15), .ZN(n_2_54));
   NOR2_X1 i_2_0_212 (.A1(n_2_0_36), .A2(n_2_0_16), .ZN(n_2_55));
   NOR2_X1 i_2_0_213 (.A1(n_2_0_36), .A2(n_2_0_17), .ZN(n_2_56));
   NOR2_X1 i_2_0_214 (.A1(n_2_0_36), .A2(n_2_0_18), .ZN(n_2_57));
   NOR2_X1 i_2_0_215 (.A1(n_2_0_36), .A2(n_2_0_19), .ZN(n_2_58));
   NOR2_X1 i_2_0_216 (.A1(n_2_0_36), .A2(n_2_0_20), .ZN(n_2_59));
   NOR2_X1 i_2_0_217 (.A1(n_2_0_36), .A2(n_2_0_21), .ZN(n_2_60));
   NOR2_X1 i_2_0_218 (.A1(n_2_0_36), .A2(n_2_0_22), .ZN(n_2_61));
   NOR2_X1 i_2_0_219 (.A1(n_2_0_36), .A2(n_2_0_23), .ZN(n_2_62));
   NOR2_X1 i_2_0_220 (.A1(n_2_0_36), .A2(n_2_0_24), .ZN(n_2_63));
   NOR2_X1 i_2_0_221 (.A1(n_2_0_36), .A2(n_2_0_25), .ZN(n_2_64));
   NOR2_X1 i_2_0_222 (.A1(n_2_0_36), .A2(n_2_0_26), .ZN(n_2_65));
   NOR2_X1 i_2_0_223 (.A1(n_2_0_36), .A2(n_2_0_27), .ZN(n_2_66));
   NOR2_X1 i_2_0_224 (.A1(n_2_0_36), .A2(n_2_0_28), .ZN(n_2_67));
   NOR2_X1 i_2_0_225 (.A1(n_2_0_36), .A2(n_2_0_29), .ZN(n_2_68));
   NOR2_X1 i_2_0_226 (.A1(n_2_0_36), .A2(n_2_0_30), .ZN(n_2_69));
   NOR2_X1 i_2_0_227 (.A1(n_2_0_36), .A2(n_2_0_31), .ZN(n_2_70));
   NOR2_X1 i_2_0_228 (.A1(n_2_0_36), .A2(n_2_0_32), .ZN(n_2_71));
   INV_X1 i_2_0_229 (.A(n_813), .ZN(n_2_0_37));
   NOR2_X1 i_2_0_230 (.A1(n_2_0_37), .A2(n_2_0_1), .ZN(n_2_72));
   NOR2_X1 i_2_0_231 (.A1(n_2_0_37), .A2(n_2_0_2), .ZN(n_2_73));
   NOR2_X1 i_2_0_232 (.A1(n_2_0_37), .A2(n_2_0_3), .ZN(n_2_74));
   NOR2_X1 i_2_0_233 (.A1(n_2_0_37), .A2(n_2_0_4), .ZN(n_2_75));
   NOR2_X1 i_2_0_234 (.A1(n_2_0_37), .A2(n_2_0_5), .ZN(n_2_76));
   NOR2_X1 i_2_0_235 (.A1(n_2_0_37), .A2(n_2_0_6), .ZN(n_2_77));
   NOR2_X1 i_2_0_236 (.A1(n_2_0_37), .A2(n_2_0_7), .ZN(n_2_78));
   NOR2_X1 i_2_0_237 (.A1(n_2_0_37), .A2(n_2_0_8), .ZN(n_2_79));
   NOR2_X1 i_2_0_238 (.A1(n_2_0_37), .A2(n_2_0_9), .ZN(n_2_80));
   NOR2_X1 i_2_0_239 (.A1(n_2_0_37), .A2(n_2_0_10), .ZN(n_2_81));
   NOR2_X1 i_2_0_240 (.A1(n_2_0_37), .A2(n_2_0_11), .ZN(n_2_82));
   NOR2_X1 i_2_0_241 (.A1(n_2_0_37), .A2(n_2_0_12), .ZN(n_2_83));
   NOR2_X1 i_2_0_242 (.A1(n_2_0_37), .A2(n_2_0_13), .ZN(n_2_84));
   NOR2_X1 i_2_0_243 (.A1(n_2_0_37), .A2(n_2_0_14), .ZN(n_2_85));
   NOR2_X1 i_2_0_244 (.A1(n_2_0_37), .A2(n_2_0_15), .ZN(n_2_86));
   NOR2_X1 i_2_0_245 (.A1(n_2_0_37), .A2(n_2_0_16), .ZN(n_2_87));
   NOR2_X1 i_2_0_246 (.A1(n_2_0_37), .A2(n_2_0_17), .ZN(n_2_88));
   NOR2_X1 i_2_0_247 (.A1(n_2_0_37), .A2(n_2_0_18), .ZN(n_2_89));
   NOR2_X1 i_2_0_248 (.A1(n_2_0_37), .A2(n_2_0_19), .ZN(n_2_90));
   NOR2_X1 i_2_0_249 (.A1(n_2_0_37), .A2(n_2_0_20), .ZN(n_2_91));
   NOR2_X1 i_2_0_250 (.A1(n_2_0_37), .A2(n_2_0_21), .ZN(n_2_92));
   NOR2_X1 i_2_0_251 (.A1(n_2_0_37), .A2(n_2_0_22), .ZN(n_2_93));
   NOR2_X1 i_2_0_252 (.A1(n_2_0_37), .A2(n_2_0_23), .ZN(n_2_94));
   NOR2_X1 i_2_0_253 (.A1(n_2_0_37), .A2(n_2_0_24), .ZN(n_2_95));
   NOR2_X1 i_2_0_254 (.A1(n_2_0_37), .A2(n_2_0_25), .ZN(n_2_96));
   NOR2_X1 i_2_0_255 (.A1(n_2_0_37), .A2(n_2_0_26), .ZN(n_2_97));
   NOR2_X1 i_2_0_256 (.A1(n_2_0_37), .A2(n_2_0_27), .ZN(n_2_98));
   NOR2_X1 i_2_0_257 (.A1(n_2_0_37), .A2(n_2_0_28), .ZN(n_2_99));
   NOR2_X1 i_2_0_258 (.A1(n_2_0_37), .A2(n_2_0_29), .ZN(n_2_100));
   NOR2_X1 i_2_0_259 (.A1(n_2_0_37), .A2(n_2_0_30), .ZN(n_2_101));
   NOR2_X1 i_2_0_260 (.A1(n_2_0_37), .A2(n_2_0_31), .ZN(n_2_102));
   NOR2_X1 i_2_0_261 (.A1(n_2_0_37), .A2(n_2_0_32), .ZN(n_2_103));
   INV_X1 i_2_0_262 (.A(n_812), .ZN(n_2_0_38));
   NOR2_X1 i_2_0_263 (.A1(n_2_0_38), .A2(n_2_0_1), .ZN(n_2_104));
   NOR2_X1 i_2_0_264 (.A1(n_2_0_38), .A2(n_2_0_2), .ZN(n_2_105));
   NOR2_X1 i_2_0_265 (.A1(n_2_0_38), .A2(n_2_0_3), .ZN(n_2_106));
   NOR2_X1 i_2_0_266 (.A1(n_2_0_38), .A2(n_2_0_4), .ZN(n_2_107));
   NOR2_X1 i_2_0_267 (.A1(n_2_0_38), .A2(n_2_0_5), .ZN(n_2_108));
   NOR2_X1 i_2_0_268 (.A1(n_2_0_38), .A2(n_2_0_6), .ZN(n_2_109));
   NOR2_X1 i_2_0_269 (.A1(n_2_0_38), .A2(n_2_0_7), .ZN(n_2_110));
   NOR2_X1 i_2_0_270 (.A1(n_2_0_38), .A2(n_2_0_8), .ZN(n_2_111));
   NOR2_X1 i_2_0_271 (.A1(n_2_0_38), .A2(n_2_0_9), .ZN(n_2_112));
   NOR2_X1 i_2_0_272 (.A1(n_2_0_38), .A2(n_2_0_10), .ZN(n_2_113));
   NOR2_X1 i_2_0_273 (.A1(n_2_0_38), .A2(n_2_0_11), .ZN(n_2_114));
   NOR2_X1 i_2_0_274 (.A1(n_2_0_38), .A2(n_2_0_12), .ZN(n_2_115));
   NOR2_X1 i_2_0_275 (.A1(n_2_0_38), .A2(n_2_0_13), .ZN(n_2_116));
   NOR2_X1 i_2_0_276 (.A1(n_2_0_38), .A2(n_2_0_14), .ZN(n_2_117));
   NOR2_X1 i_2_0_277 (.A1(n_2_0_38), .A2(n_2_0_15), .ZN(n_2_118));
   NOR2_X1 i_2_0_278 (.A1(n_2_0_38), .A2(n_2_0_16), .ZN(n_2_119));
   NOR2_X1 i_2_0_279 (.A1(n_2_0_38), .A2(n_2_0_17), .ZN(n_2_120));
   NOR2_X1 i_2_0_280 (.A1(n_2_0_38), .A2(n_2_0_18), .ZN(n_2_121));
   NOR2_X1 i_2_0_281 (.A1(n_2_0_38), .A2(n_2_0_19), .ZN(n_2_122));
   NOR2_X1 i_2_0_282 (.A1(n_2_0_38), .A2(n_2_0_20), .ZN(n_2_123));
   NOR2_X1 i_2_0_283 (.A1(n_2_0_38), .A2(n_2_0_21), .ZN(n_2_124));
   NOR2_X1 i_2_0_284 (.A1(n_2_0_38), .A2(n_2_0_22), .ZN(n_2_125));
   NOR2_X1 i_2_0_285 (.A1(n_2_0_38), .A2(n_2_0_23), .ZN(n_2_126));
   NOR2_X1 i_2_0_286 (.A1(n_2_0_38), .A2(n_2_0_24), .ZN(n_2_127));
   NOR2_X1 i_2_0_287 (.A1(n_2_0_38), .A2(n_2_0_25), .ZN(n_2_128));
   NOR2_X1 i_2_0_288 (.A1(n_2_0_38), .A2(n_2_0_26), .ZN(n_2_129));
   NOR2_X1 i_2_0_289 (.A1(n_2_0_38), .A2(n_2_0_27), .ZN(n_2_130));
   NOR2_X1 i_2_0_290 (.A1(n_2_0_38), .A2(n_2_0_28), .ZN(n_2_131));
   NOR2_X1 i_2_0_291 (.A1(n_2_0_38), .A2(n_2_0_29), .ZN(n_2_132));
   NOR2_X1 i_2_0_292 (.A1(n_2_0_38), .A2(n_2_0_30), .ZN(n_2_133));
   NOR2_X1 i_2_0_293 (.A1(n_2_0_38), .A2(n_2_0_31), .ZN(n_2_134));
   NOR2_X1 i_2_0_294 (.A1(n_2_0_38), .A2(n_2_0_32), .ZN(n_2_135));
   INV_X1 i_2_0_295 (.A(n_811), .ZN(n_2_0_39));
   NOR2_X1 i_2_0_296 (.A1(n_2_0_39), .A2(n_2_0_1), .ZN(n_161));
   NOR2_X1 i_2_0_297 (.A1(n_2_0_39), .A2(n_2_0_2), .ZN(n_2_136));
   NOR2_X1 i_2_0_298 (.A1(n_2_0_39), .A2(n_2_0_3), .ZN(n_2_137));
   NOR2_X1 i_2_0_299 (.A1(n_2_0_39), .A2(n_2_0_4), .ZN(n_2_138));
   NOR2_X1 i_2_0_300 (.A1(n_2_0_39), .A2(n_2_0_5), .ZN(n_2_139));
   NOR2_X1 i_2_0_301 (.A1(n_2_0_39), .A2(n_2_0_6), .ZN(n_2_140));
   NOR2_X1 i_2_0_302 (.A1(n_2_0_39), .A2(n_2_0_7), .ZN(n_2_141));
   NOR2_X1 i_2_0_303 (.A1(n_2_0_39), .A2(n_2_0_8), .ZN(n_2_142));
   NOR2_X1 i_2_0_304 (.A1(n_2_0_39), .A2(n_2_0_9), .ZN(n_2_143));
   NOR2_X1 i_2_0_305 (.A1(n_2_0_39), .A2(n_2_0_10), .ZN(n_2_144));
   NOR2_X1 i_2_0_306 (.A1(n_2_0_39), .A2(n_2_0_11), .ZN(n_2_145));
   NOR2_X1 i_2_0_307 (.A1(n_2_0_39), .A2(n_2_0_12), .ZN(n_2_146));
   NOR2_X1 i_2_0_308 (.A1(n_2_0_39), .A2(n_2_0_13), .ZN(n_2_147));
   NOR2_X1 i_2_0_309 (.A1(n_2_0_39), .A2(n_2_0_14), .ZN(n_2_148));
   NOR2_X1 i_2_0_310 (.A1(n_2_0_39), .A2(n_2_0_15), .ZN(n_2_149));
   NOR2_X1 i_2_0_311 (.A1(n_2_0_39), .A2(n_2_0_16), .ZN(n_2_150));
   NOR2_X1 i_2_0_312 (.A1(n_2_0_39), .A2(n_2_0_17), .ZN(n_2_151));
   NOR2_X1 i_2_0_313 (.A1(n_2_0_39), .A2(n_2_0_18), .ZN(n_2_152));
   NOR2_X1 i_2_0_314 (.A1(n_2_0_39), .A2(n_2_0_19), .ZN(n_2_153));
   NOR2_X1 i_2_0_315 (.A1(n_2_0_39), .A2(n_2_0_20), .ZN(n_2_154));
   NOR2_X1 i_2_0_316 (.A1(n_2_0_39), .A2(n_2_0_21), .ZN(n_2_155));
   NOR2_X1 i_2_0_317 (.A1(n_2_0_39), .A2(n_2_0_22), .ZN(n_2_156));
   NOR2_X1 i_2_0_318 (.A1(n_2_0_39), .A2(n_2_0_23), .ZN(n_2_157));
   NOR2_X1 i_2_0_319 (.A1(n_2_0_39), .A2(n_2_0_24), .ZN(n_2_158));
   NOR2_X1 i_2_0_320 (.A1(n_2_0_39), .A2(n_2_0_25), .ZN(n_2_159));
   NOR2_X1 i_2_0_321 (.A1(n_2_0_39), .A2(n_2_0_26), .ZN(n_2_160));
   NOR2_X1 i_2_0_322 (.A1(n_2_0_39), .A2(n_2_0_27), .ZN(n_2_161));
   NOR2_X1 i_2_0_323 (.A1(n_2_0_39), .A2(n_2_0_28), .ZN(n_2_162));
   NOR2_X1 i_2_0_324 (.A1(n_2_0_39), .A2(n_2_0_29), .ZN(n_2_163));
   NOR2_X1 i_2_0_325 (.A1(n_2_0_39), .A2(n_2_0_30), .ZN(n_2_164));
   NOR2_X1 i_2_0_326 (.A1(n_2_0_39), .A2(n_2_0_31), .ZN(n_2_165));
   NOR2_X1 i_2_0_327 (.A1(n_2_0_39), .A2(n_2_0_32), .ZN(n_2_166));
   INV_X1 i_2_0_328 (.A(n_810), .ZN(n_2_0_40));
   NOR2_X1 i_2_0_329 (.A1(n_2_0_40), .A2(n_2_0_1), .ZN(n_2_167));
   NOR2_X1 i_2_0_330 (.A1(n_2_0_40), .A2(n_2_0_2), .ZN(n_2_168));
   NOR2_X1 i_2_0_331 (.A1(n_2_0_40), .A2(n_2_0_3), .ZN(n_2_169));
   NOR2_X1 i_2_0_332 (.A1(n_2_0_40), .A2(n_2_0_4), .ZN(n_2_170));
   NOR2_X1 i_2_0_333 (.A1(n_2_0_40), .A2(n_2_0_5), .ZN(n_2_171));
   NOR2_X1 i_2_0_334 (.A1(n_2_0_40), .A2(n_2_0_6), .ZN(n_2_172));
   NOR2_X1 i_2_0_335 (.A1(n_2_0_40), .A2(n_2_0_7), .ZN(n_2_173));
   NOR2_X1 i_2_0_336 (.A1(n_2_0_40), .A2(n_2_0_8), .ZN(n_2_174));
   NOR2_X1 i_2_0_337 (.A1(n_2_0_40), .A2(n_2_0_9), .ZN(n_2_175));
   NOR2_X1 i_2_0_338 (.A1(n_2_0_40), .A2(n_2_0_10), .ZN(n_2_176));
   NOR2_X1 i_2_0_339 (.A1(n_2_0_40), .A2(n_2_0_11), .ZN(n_2_177));
   NOR2_X1 i_2_0_340 (.A1(n_2_0_40), .A2(n_2_0_12), .ZN(n_2_178));
   NOR2_X1 i_2_0_341 (.A1(n_2_0_40), .A2(n_2_0_13), .ZN(n_2_179));
   NOR2_X1 i_2_0_342 (.A1(n_2_0_40), .A2(n_2_0_14), .ZN(n_2_180));
   NOR2_X1 i_2_0_343 (.A1(n_2_0_40), .A2(n_2_0_15), .ZN(n_2_181));
   NOR2_X1 i_2_0_344 (.A1(n_2_0_40), .A2(n_2_0_16), .ZN(n_2_182));
   NOR2_X1 i_2_0_345 (.A1(n_2_0_40), .A2(n_2_0_17), .ZN(n_2_183));
   NOR2_X1 i_2_0_346 (.A1(n_2_0_40), .A2(n_2_0_18), .ZN(n_2_184));
   NOR2_X1 i_2_0_347 (.A1(n_2_0_40), .A2(n_2_0_19), .ZN(n_2_185));
   NOR2_X1 i_2_0_348 (.A1(n_2_0_40), .A2(n_2_0_20), .ZN(n_2_186));
   NOR2_X1 i_2_0_349 (.A1(n_2_0_40), .A2(n_2_0_21), .ZN(n_2_187));
   NOR2_X1 i_2_0_350 (.A1(n_2_0_40), .A2(n_2_0_22), .ZN(n_2_188));
   NOR2_X1 i_2_0_351 (.A1(n_2_0_40), .A2(n_2_0_23), .ZN(n_2_189));
   NOR2_X1 i_2_0_352 (.A1(n_2_0_40), .A2(n_2_0_24), .ZN(n_2_190));
   NOR2_X1 i_2_0_353 (.A1(n_2_0_40), .A2(n_2_0_25), .ZN(n_2_191));
   NOR2_X1 i_2_0_354 (.A1(n_2_0_40), .A2(n_2_0_26), .ZN(n_2_192));
   NOR2_X1 i_2_0_355 (.A1(n_2_0_40), .A2(n_2_0_27), .ZN(n_2_193));
   NOR2_X1 i_2_0_356 (.A1(n_2_0_40), .A2(n_2_0_28), .ZN(n_2_194));
   NOR2_X1 i_2_0_357 (.A1(n_2_0_40), .A2(n_2_0_29), .ZN(n_2_195));
   NOR2_X1 i_2_0_358 (.A1(n_2_0_40), .A2(n_2_0_30), .ZN(n_2_196));
   NOR2_X1 i_2_0_359 (.A1(n_2_0_40), .A2(n_2_0_31), .ZN(n_2_197));
   NOR2_X1 i_2_0_360 (.A1(n_2_0_40), .A2(n_2_0_32), .ZN(n_2_198));
   INV_X1 i_2_0_361 (.A(n_809), .ZN(n_2_0_41));
   NOR2_X1 i_2_0_362 (.A1(n_2_0_41), .A2(n_2_0_1), .ZN(n_2_199));
   NOR2_X1 i_2_0_363 (.A1(n_2_0_41), .A2(n_2_0_2), .ZN(n_2_200));
   NOR2_X1 i_2_0_364 (.A1(n_2_0_41), .A2(n_2_0_3), .ZN(n_2_201));
   NOR2_X1 i_2_0_365 (.A1(n_2_0_41), .A2(n_2_0_4), .ZN(n_2_202));
   NOR2_X1 i_2_0_366 (.A1(n_2_0_41), .A2(n_2_0_5), .ZN(n_2_203));
   NOR2_X1 i_2_0_367 (.A1(n_2_0_41), .A2(n_2_0_6), .ZN(n_2_204));
   NOR2_X1 i_2_0_368 (.A1(n_2_0_41), .A2(n_2_0_7), .ZN(n_2_205));
   NOR2_X1 i_2_0_369 (.A1(n_2_0_41), .A2(n_2_0_8), .ZN(n_2_206));
   NOR2_X1 i_2_0_370 (.A1(n_2_0_41), .A2(n_2_0_9), .ZN(n_2_207));
   NOR2_X1 i_2_0_371 (.A1(n_2_0_41), .A2(n_2_0_10), .ZN(n_2_208));
   NOR2_X1 i_2_0_372 (.A1(n_2_0_41), .A2(n_2_0_11), .ZN(n_2_209));
   NOR2_X1 i_2_0_373 (.A1(n_2_0_41), .A2(n_2_0_12), .ZN(n_2_210));
   NOR2_X1 i_2_0_374 (.A1(n_2_0_41), .A2(n_2_0_13), .ZN(n_2_211));
   NOR2_X1 i_2_0_375 (.A1(n_2_0_41), .A2(n_2_0_14), .ZN(n_2_212));
   NOR2_X1 i_2_0_376 (.A1(n_2_0_41), .A2(n_2_0_15), .ZN(n_2_213));
   NOR2_X1 i_2_0_377 (.A1(n_2_0_41), .A2(n_2_0_16), .ZN(n_2_214));
   NOR2_X1 i_2_0_378 (.A1(n_2_0_41), .A2(n_2_0_17), .ZN(n_2_215));
   NOR2_X1 i_2_0_379 (.A1(n_2_0_41), .A2(n_2_0_18), .ZN(n_2_216));
   NOR2_X1 i_2_0_380 (.A1(n_2_0_41), .A2(n_2_0_19), .ZN(n_2_217));
   NOR2_X1 i_2_0_381 (.A1(n_2_0_41), .A2(n_2_0_20), .ZN(n_2_218));
   NOR2_X1 i_2_0_382 (.A1(n_2_0_41), .A2(n_2_0_21), .ZN(n_2_219));
   NOR2_X1 i_2_0_383 (.A1(n_2_0_41), .A2(n_2_0_22), .ZN(n_2_220));
   NOR2_X1 i_2_0_384 (.A1(n_2_0_41), .A2(n_2_0_23), .ZN(n_2_221));
   NOR2_X1 i_2_0_385 (.A1(n_2_0_41), .A2(n_2_0_24), .ZN(n_2_222));
   NOR2_X1 i_2_0_386 (.A1(n_2_0_41), .A2(n_2_0_25), .ZN(n_2_223));
   NOR2_X1 i_2_0_387 (.A1(n_2_0_41), .A2(n_2_0_26), .ZN(n_2_224));
   NOR2_X1 i_2_0_388 (.A1(n_2_0_41), .A2(n_2_0_27), .ZN(n_2_225));
   NOR2_X1 i_2_0_389 (.A1(n_2_0_41), .A2(n_2_0_28), .ZN(n_2_226));
   NOR2_X1 i_2_0_390 (.A1(n_2_0_41), .A2(n_2_0_29), .ZN(n_2_227));
   NOR2_X1 i_2_0_391 (.A1(n_2_0_41), .A2(n_2_0_30), .ZN(n_2_228));
   NOR2_X1 i_2_0_392 (.A1(n_2_0_41), .A2(n_2_0_31), .ZN(n_2_229));
   NOR2_X1 i_2_0_393 (.A1(n_2_0_41), .A2(n_2_0_32), .ZN(n_2_230));
   INV_X1 i_2_0_394 (.A(n_808), .ZN(n_2_0_42));
   NOR2_X1 i_2_0_395 (.A1(n_2_0_42), .A2(n_2_0_1), .ZN(n_162));
   NOR2_X1 i_2_0_396 (.A1(n_2_0_42), .A2(n_2_0_2), .ZN(n_2_231));
   NOR2_X1 i_2_0_397 (.A1(n_2_0_42), .A2(n_2_0_3), .ZN(n_2_232));
   NOR2_X1 i_2_0_398 (.A1(n_2_0_42), .A2(n_2_0_4), .ZN(n_2_233));
   NOR2_X1 i_2_0_399 (.A1(n_2_0_42), .A2(n_2_0_5), .ZN(n_2_234));
   NOR2_X1 i_2_0_400 (.A1(n_2_0_42), .A2(n_2_0_6), .ZN(n_2_235));
   NOR2_X1 i_2_0_401 (.A1(n_2_0_42), .A2(n_2_0_7), .ZN(n_2_236));
   NOR2_X1 i_2_0_402 (.A1(n_2_0_42), .A2(n_2_0_8), .ZN(n_2_237));
   NOR2_X1 i_2_0_403 (.A1(n_2_0_42), .A2(n_2_0_9), .ZN(n_2_238));
   NOR2_X1 i_2_0_404 (.A1(n_2_0_42), .A2(n_2_0_10), .ZN(n_2_239));
   NOR2_X1 i_2_0_405 (.A1(n_2_0_42), .A2(n_2_0_11), .ZN(n_2_240));
   NOR2_X1 i_2_0_406 (.A1(n_2_0_42), .A2(n_2_0_12), .ZN(n_2_241));
   NOR2_X1 i_2_0_407 (.A1(n_2_0_42), .A2(n_2_0_13), .ZN(n_2_242));
   NOR2_X1 i_2_0_408 (.A1(n_2_0_42), .A2(n_2_0_14), .ZN(n_2_243));
   NOR2_X1 i_2_0_409 (.A1(n_2_0_42), .A2(n_2_0_15), .ZN(n_2_244));
   NOR2_X1 i_2_0_410 (.A1(n_2_0_42), .A2(n_2_0_16), .ZN(n_2_245));
   NOR2_X1 i_2_0_411 (.A1(n_2_0_42), .A2(n_2_0_17), .ZN(n_2_246));
   NOR2_X1 i_2_0_412 (.A1(n_2_0_42), .A2(n_2_0_18), .ZN(n_2_247));
   NOR2_X1 i_2_0_413 (.A1(n_2_0_42), .A2(n_2_0_19), .ZN(n_2_248));
   NOR2_X1 i_2_0_414 (.A1(n_2_0_42), .A2(n_2_0_20), .ZN(n_2_249));
   NOR2_X1 i_2_0_415 (.A1(n_2_0_42), .A2(n_2_0_21), .ZN(n_2_250));
   NOR2_X1 i_2_0_416 (.A1(n_2_0_42), .A2(n_2_0_22), .ZN(n_2_251));
   NOR2_X1 i_2_0_417 (.A1(n_2_0_42), .A2(n_2_0_23), .ZN(n_2_252));
   NOR2_X1 i_2_0_418 (.A1(n_2_0_42), .A2(n_2_0_24), .ZN(n_2_253));
   NOR2_X1 i_2_0_419 (.A1(n_2_0_42), .A2(n_2_0_25), .ZN(n_2_254));
   NOR2_X1 i_2_0_420 (.A1(n_2_0_42), .A2(n_2_0_26), .ZN(n_2_255));
   NOR2_X1 i_2_0_421 (.A1(n_2_0_42), .A2(n_2_0_27), .ZN(n_2_256));
   NOR2_X1 i_2_0_422 (.A1(n_2_0_42), .A2(n_2_0_28), .ZN(n_2_257));
   NOR2_X1 i_2_0_423 (.A1(n_2_0_42), .A2(n_2_0_29), .ZN(n_2_258));
   NOR2_X1 i_2_0_424 (.A1(n_2_0_42), .A2(n_2_0_30), .ZN(n_2_259));
   NOR2_X1 i_2_0_425 (.A1(n_2_0_42), .A2(n_2_0_31), .ZN(n_2_260));
   NOR2_X1 i_2_0_426 (.A1(n_2_0_42), .A2(n_2_0_32), .ZN(n_2_261));
   INV_X1 i_2_0_427 (.A(n_807), .ZN(n_2_0_43));
   NOR2_X1 i_2_0_428 (.A1(n_2_0_43), .A2(n_2_0_1), .ZN(n_2_262));
   NOR2_X1 i_2_0_429 (.A1(n_2_0_43), .A2(n_2_0_2), .ZN(n_2_263));
   NOR2_X1 i_2_0_430 (.A1(n_2_0_43), .A2(n_2_0_3), .ZN(n_2_264));
   NOR2_X1 i_2_0_431 (.A1(n_2_0_43), .A2(n_2_0_4), .ZN(n_2_265));
   NOR2_X1 i_2_0_432 (.A1(n_2_0_43), .A2(n_2_0_5), .ZN(n_2_266));
   NOR2_X1 i_2_0_433 (.A1(n_2_0_43), .A2(n_2_0_6), .ZN(n_2_267));
   NOR2_X1 i_2_0_434 (.A1(n_2_0_43), .A2(n_2_0_7), .ZN(n_2_268));
   NOR2_X1 i_2_0_435 (.A1(n_2_0_43), .A2(n_2_0_8), .ZN(n_2_269));
   NOR2_X1 i_2_0_436 (.A1(n_2_0_43), .A2(n_2_0_9), .ZN(n_2_270));
   NOR2_X1 i_2_0_437 (.A1(n_2_0_43), .A2(n_2_0_10), .ZN(n_2_271));
   NOR2_X1 i_2_0_438 (.A1(n_2_0_43), .A2(n_2_0_11), .ZN(n_2_272));
   NOR2_X1 i_2_0_439 (.A1(n_2_0_43), .A2(n_2_0_12), .ZN(n_2_273));
   NOR2_X1 i_2_0_440 (.A1(n_2_0_43), .A2(n_2_0_13), .ZN(n_2_274));
   NOR2_X1 i_2_0_441 (.A1(n_2_0_43), .A2(n_2_0_14), .ZN(n_2_275));
   NOR2_X1 i_2_0_442 (.A1(n_2_0_43), .A2(n_2_0_15), .ZN(n_2_276));
   NOR2_X1 i_2_0_443 (.A1(n_2_0_43), .A2(n_2_0_16), .ZN(n_2_277));
   NOR2_X1 i_2_0_444 (.A1(n_2_0_43), .A2(n_2_0_17), .ZN(n_2_278));
   NOR2_X1 i_2_0_445 (.A1(n_2_0_43), .A2(n_2_0_18), .ZN(n_2_279));
   NOR2_X1 i_2_0_446 (.A1(n_2_0_43), .A2(n_2_0_19), .ZN(n_2_280));
   NOR2_X1 i_2_0_447 (.A1(n_2_0_43), .A2(n_2_0_20), .ZN(n_2_281));
   NOR2_X1 i_2_0_448 (.A1(n_2_0_43), .A2(n_2_0_21), .ZN(n_2_282));
   NOR2_X1 i_2_0_449 (.A1(n_2_0_43), .A2(n_2_0_22), .ZN(n_2_283));
   NOR2_X1 i_2_0_450 (.A1(n_2_0_43), .A2(n_2_0_23), .ZN(n_2_284));
   NOR2_X1 i_2_0_451 (.A1(n_2_0_43), .A2(n_2_0_24), .ZN(n_2_285));
   NOR2_X1 i_2_0_452 (.A1(n_2_0_43), .A2(n_2_0_25), .ZN(n_2_286));
   NOR2_X1 i_2_0_453 (.A1(n_2_0_43), .A2(n_2_0_26), .ZN(n_2_287));
   NOR2_X1 i_2_0_454 (.A1(n_2_0_43), .A2(n_2_0_27), .ZN(n_2_288));
   NOR2_X1 i_2_0_455 (.A1(n_2_0_43), .A2(n_2_0_28), .ZN(n_2_289));
   NOR2_X1 i_2_0_456 (.A1(n_2_0_43), .A2(n_2_0_29), .ZN(n_2_290));
   NOR2_X1 i_2_0_457 (.A1(n_2_0_43), .A2(n_2_0_30), .ZN(n_2_291));
   NOR2_X1 i_2_0_458 (.A1(n_2_0_43), .A2(n_2_0_31), .ZN(n_2_292));
   NOR2_X1 i_2_0_459 (.A1(n_2_0_43), .A2(n_2_0_32), .ZN(n_2_293));
   INV_X1 i_2_0_460 (.A(n_806), .ZN(n_2_0_44));
   NOR2_X1 i_2_0_461 (.A1(n_2_0_44), .A2(n_2_0_1), .ZN(n_2_294));
   NOR2_X1 i_2_0_462 (.A1(n_2_0_44), .A2(n_2_0_2), .ZN(n_2_295));
   NOR2_X1 i_2_0_463 (.A1(n_2_0_44), .A2(n_2_0_3), .ZN(n_2_296));
   NOR2_X1 i_2_0_464 (.A1(n_2_0_44), .A2(n_2_0_4), .ZN(n_2_297));
   NOR2_X1 i_2_0_465 (.A1(n_2_0_44), .A2(n_2_0_5), .ZN(n_2_298));
   NOR2_X1 i_2_0_466 (.A1(n_2_0_44), .A2(n_2_0_6), .ZN(n_2_299));
   NOR2_X1 i_2_0_467 (.A1(n_2_0_44), .A2(n_2_0_7), .ZN(n_2_300));
   NOR2_X1 i_2_0_468 (.A1(n_2_0_44), .A2(n_2_0_8), .ZN(n_2_301));
   NOR2_X1 i_2_0_469 (.A1(n_2_0_44), .A2(n_2_0_9), .ZN(n_2_302));
   NOR2_X1 i_2_0_470 (.A1(n_2_0_44), .A2(n_2_0_10), .ZN(n_2_303));
   NOR2_X1 i_2_0_471 (.A1(n_2_0_44), .A2(n_2_0_11), .ZN(n_2_304));
   NOR2_X1 i_2_0_472 (.A1(n_2_0_44), .A2(n_2_0_12), .ZN(n_2_305));
   NOR2_X1 i_2_0_473 (.A1(n_2_0_44), .A2(n_2_0_13), .ZN(n_2_306));
   NOR2_X1 i_2_0_474 (.A1(n_2_0_44), .A2(n_2_0_14), .ZN(n_2_307));
   NOR2_X1 i_2_0_475 (.A1(n_2_0_44), .A2(n_2_0_15), .ZN(n_2_308));
   NOR2_X1 i_2_0_476 (.A1(n_2_0_44), .A2(n_2_0_16), .ZN(n_2_309));
   NOR2_X1 i_2_0_477 (.A1(n_2_0_44), .A2(n_2_0_17), .ZN(n_2_310));
   NOR2_X1 i_2_0_478 (.A1(n_2_0_44), .A2(n_2_0_18), .ZN(n_2_311));
   NOR2_X1 i_2_0_479 (.A1(n_2_0_44), .A2(n_2_0_19), .ZN(n_2_312));
   NOR2_X1 i_2_0_480 (.A1(n_2_0_44), .A2(n_2_0_20), .ZN(n_2_313));
   NOR2_X1 i_2_0_481 (.A1(n_2_0_44), .A2(n_2_0_21), .ZN(n_2_314));
   NOR2_X1 i_2_0_482 (.A1(n_2_0_44), .A2(n_2_0_22), .ZN(n_2_315));
   NOR2_X1 i_2_0_483 (.A1(n_2_0_44), .A2(n_2_0_23), .ZN(n_2_316));
   NOR2_X1 i_2_0_484 (.A1(n_2_0_44), .A2(n_2_0_24), .ZN(n_2_317));
   NOR2_X1 i_2_0_485 (.A1(n_2_0_44), .A2(n_2_0_25), .ZN(n_2_318));
   NOR2_X1 i_2_0_486 (.A1(n_2_0_44), .A2(n_2_0_26), .ZN(n_2_319));
   NOR2_X1 i_2_0_487 (.A1(n_2_0_44), .A2(n_2_0_27), .ZN(n_2_320));
   NOR2_X1 i_2_0_488 (.A1(n_2_0_44), .A2(n_2_0_28), .ZN(n_2_321));
   NOR2_X1 i_2_0_489 (.A1(n_2_0_44), .A2(n_2_0_29), .ZN(n_2_322));
   NOR2_X1 i_2_0_490 (.A1(n_2_0_44), .A2(n_2_0_30), .ZN(n_2_323));
   NOR2_X1 i_2_0_491 (.A1(n_2_0_44), .A2(n_2_0_31), .ZN(n_2_324));
   NOR2_X1 i_2_0_492 (.A1(n_2_0_44), .A2(n_2_0_32), .ZN(n_2_325));
   INV_X1 i_2_0_493 (.A(n_805), .ZN(n_2_0_45));
   NOR2_X1 i_2_0_494 (.A1(n_2_0_45), .A2(n_2_0_1), .ZN(n_163));
   NOR2_X1 i_2_0_495 (.A1(n_2_0_45), .A2(n_2_0_2), .ZN(n_2_326));
   NOR2_X1 i_2_0_496 (.A1(n_2_0_45), .A2(n_2_0_3), .ZN(n_2_327));
   NOR2_X1 i_2_0_497 (.A1(n_2_0_45), .A2(n_2_0_4), .ZN(n_2_328));
   NOR2_X1 i_2_0_498 (.A1(n_2_0_45), .A2(n_2_0_5), .ZN(n_2_329));
   NOR2_X1 i_2_0_499 (.A1(n_2_0_45), .A2(n_2_0_6), .ZN(n_2_330));
   NOR2_X1 i_2_0_500 (.A1(n_2_0_45), .A2(n_2_0_7), .ZN(n_2_331));
   NOR2_X1 i_2_0_501 (.A1(n_2_0_45), .A2(n_2_0_8), .ZN(n_2_332));
   NOR2_X1 i_2_0_502 (.A1(n_2_0_45), .A2(n_2_0_9), .ZN(n_2_333));
   NOR2_X1 i_2_0_503 (.A1(n_2_0_45), .A2(n_2_0_10), .ZN(n_2_334));
   NOR2_X1 i_2_0_504 (.A1(n_2_0_45), .A2(n_2_0_11), .ZN(n_2_335));
   NOR2_X1 i_2_0_505 (.A1(n_2_0_45), .A2(n_2_0_12), .ZN(n_2_336));
   NOR2_X1 i_2_0_506 (.A1(n_2_0_45), .A2(n_2_0_13), .ZN(n_2_337));
   NOR2_X1 i_2_0_507 (.A1(n_2_0_45), .A2(n_2_0_14), .ZN(n_2_338));
   NOR2_X1 i_2_0_508 (.A1(n_2_0_45), .A2(n_2_0_15), .ZN(n_2_339));
   NOR2_X1 i_2_0_509 (.A1(n_2_0_45), .A2(n_2_0_16), .ZN(n_2_340));
   NOR2_X1 i_2_0_510 (.A1(n_2_0_45), .A2(n_2_0_17), .ZN(n_2_341));
   NOR2_X1 i_2_0_511 (.A1(n_2_0_45), .A2(n_2_0_18), .ZN(n_2_342));
   NOR2_X1 i_2_0_512 (.A1(n_2_0_45), .A2(n_2_0_19), .ZN(n_2_343));
   NOR2_X1 i_2_0_513 (.A1(n_2_0_45), .A2(n_2_0_20), .ZN(n_2_344));
   NOR2_X1 i_2_0_514 (.A1(n_2_0_45), .A2(n_2_0_21), .ZN(n_2_345));
   NOR2_X1 i_2_0_515 (.A1(n_2_0_45), .A2(n_2_0_22), .ZN(n_2_346));
   NOR2_X1 i_2_0_516 (.A1(n_2_0_45), .A2(n_2_0_23), .ZN(n_2_347));
   NOR2_X1 i_2_0_517 (.A1(n_2_0_45), .A2(n_2_0_24), .ZN(n_2_348));
   NOR2_X1 i_2_0_518 (.A1(n_2_0_45), .A2(n_2_0_25), .ZN(n_2_349));
   NOR2_X1 i_2_0_519 (.A1(n_2_0_45), .A2(n_2_0_26), .ZN(n_2_350));
   NOR2_X1 i_2_0_520 (.A1(n_2_0_45), .A2(n_2_0_27), .ZN(n_2_351));
   NOR2_X1 i_2_0_521 (.A1(n_2_0_45), .A2(n_2_0_28), .ZN(n_2_352));
   NOR2_X1 i_2_0_522 (.A1(n_2_0_45), .A2(n_2_0_29), .ZN(n_2_353));
   NOR2_X1 i_2_0_523 (.A1(n_2_0_45), .A2(n_2_0_30), .ZN(n_2_354));
   NOR2_X1 i_2_0_524 (.A1(n_2_0_45), .A2(n_2_0_31), .ZN(n_2_355));
   NOR2_X1 i_2_0_525 (.A1(n_2_0_45), .A2(n_2_0_32), .ZN(n_2_356));
   INV_X1 i_2_0_526 (.A(n_804), .ZN(n_2_0_46));
   NOR2_X1 i_2_0_527 (.A1(n_2_0_46), .A2(n_2_0_1), .ZN(n_2_357));
   NOR2_X1 i_2_0_528 (.A1(n_2_0_46), .A2(n_2_0_2), .ZN(n_2_358));
   NOR2_X1 i_2_0_529 (.A1(n_2_0_46), .A2(n_2_0_3), .ZN(n_2_359));
   NOR2_X1 i_2_0_530 (.A1(n_2_0_46), .A2(n_2_0_4), .ZN(n_2_360));
   NOR2_X1 i_2_0_531 (.A1(n_2_0_46), .A2(n_2_0_5), .ZN(n_2_361));
   NOR2_X1 i_2_0_532 (.A1(n_2_0_46), .A2(n_2_0_6), .ZN(n_2_362));
   NOR2_X1 i_2_0_533 (.A1(n_2_0_46), .A2(n_2_0_7), .ZN(n_2_363));
   NOR2_X1 i_2_0_534 (.A1(n_2_0_46), .A2(n_2_0_8), .ZN(n_2_364));
   NOR2_X1 i_2_0_535 (.A1(n_2_0_46), .A2(n_2_0_9), .ZN(n_2_365));
   NOR2_X1 i_2_0_536 (.A1(n_2_0_46), .A2(n_2_0_10), .ZN(n_2_366));
   NOR2_X1 i_2_0_537 (.A1(n_2_0_46), .A2(n_2_0_11), .ZN(n_2_367));
   NOR2_X1 i_2_0_538 (.A1(n_2_0_46), .A2(n_2_0_12), .ZN(n_2_368));
   NOR2_X1 i_2_0_539 (.A1(n_2_0_46), .A2(n_2_0_13), .ZN(n_2_369));
   NOR2_X1 i_2_0_540 (.A1(n_2_0_46), .A2(n_2_0_14), .ZN(n_2_370));
   NOR2_X1 i_2_0_541 (.A1(n_2_0_46), .A2(n_2_0_15), .ZN(n_2_371));
   NOR2_X1 i_2_0_542 (.A1(n_2_0_46), .A2(n_2_0_16), .ZN(n_2_372));
   NOR2_X1 i_2_0_543 (.A1(n_2_0_46), .A2(n_2_0_17), .ZN(n_2_373));
   NOR2_X1 i_2_0_544 (.A1(n_2_0_46), .A2(n_2_0_18), .ZN(n_2_374));
   NOR2_X1 i_2_0_545 (.A1(n_2_0_46), .A2(n_2_0_19), .ZN(n_2_375));
   NOR2_X1 i_2_0_546 (.A1(n_2_0_46), .A2(n_2_0_20), .ZN(n_2_376));
   NOR2_X1 i_2_0_547 (.A1(n_2_0_46), .A2(n_2_0_21), .ZN(n_2_377));
   NOR2_X1 i_2_0_548 (.A1(n_2_0_46), .A2(n_2_0_22), .ZN(n_2_378));
   NOR2_X1 i_2_0_549 (.A1(n_2_0_46), .A2(n_2_0_23), .ZN(n_2_379));
   NOR2_X1 i_2_0_550 (.A1(n_2_0_46), .A2(n_2_0_24), .ZN(n_2_380));
   NOR2_X1 i_2_0_551 (.A1(n_2_0_46), .A2(n_2_0_25), .ZN(n_2_381));
   NOR2_X1 i_2_0_552 (.A1(n_2_0_46), .A2(n_2_0_26), .ZN(n_2_382));
   NOR2_X1 i_2_0_553 (.A1(n_2_0_46), .A2(n_2_0_27), .ZN(n_2_383));
   NOR2_X1 i_2_0_554 (.A1(n_2_0_46), .A2(n_2_0_28), .ZN(n_2_384));
   NOR2_X1 i_2_0_555 (.A1(n_2_0_46), .A2(n_2_0_29), .ZN(n_2_385));
   NOR2_X1 i_2_0_556 (.A1(n_2_0_46), .A2(n_2_0_30), .ZN(n_2_386));
   NOR2_X1 i_2_0_557 (.A1(n_2_0_46), .A2(n_2_0_31), .ZN(n_2_387));
   NOR2_X1 i_2_0_558 (.A1(n_2_0_46), .A2(n_2_0_32), .ZN(n_2_388));
   INV_X1 i_2_0_559 (.A(n_803), .ZN(n_2_0_47));
   NOR2_X1 i_2_0_560 (.A1(n_2_0_47), .A2(n_2_0_1), .ZN(n_2_389));
   NOR2_X1 i_2_0_561 (.A1(n_2_0_47), .A2(n_2_0_2), .ZN(n_2_390));
   NOR2_X1 i_2_0_562 (.A1(n_2_0_47), .A2(n_2_0_3), .ZN(n_2_391));
   NOR2_X1 i_2_0_563 (.A1(n_2_0_47), .A2(n_2_0_4), .ZN(n_2_392));
   NOR2_X1 i_2_0_564 (.A1(n_2_0_47), .A2(n_2_0_5), .ZN(n_2_393));
   NOR2_X1 i_2_0_565 (.A1(n_2_0_47), .A2(n_2_0_6), .ZN(n_2_394));
   NOR2_X1 i_2_0_566 (.A1(n_2_0_47), .A2(n_2_0_7), .ZN(n_2_395));
   NOR2_X1 i_2_0_567 (.A1(n_2_0_47), .A2(n_2_0_8), .ZN(n_2_396));
   NOR2_X1 i_2_0_568 (.A1(n_2_0_47), .A2(n_2_0_9), .ZN(n_2_397));
   NOR2_X1 i_2_0_569 (.A1(n_2_0_47), .A2(n_2_0_10), .ZN(n_2_398));
   NOR2_X1 i_2_0_570 (.A1(n_2_0_47), .A2(n_2_0_11), .ZN(n_2_399));
   NOR2_X1 i_2_0_571 (.A1(n_2_0_47), .A2(n_2_0_12), .ZN(n_2_400));
   NOR2_X1 i_2_0_572 (.A1(n_2_0_47), .A2(n_2_0_13), .ZN(n_2_401));
   NOR2_X1 i_2_0_573 (.A1(n_2_0_47), .A2(n_2_0_14), .ZN(n_2_402));
   NOR2_X1 i_2_0_574 (.A1(n_2_0_47), .A2(n_2_0_15), .ZN(n_2_403));
   NOR2_X1 i_2_0_575 (.A1(n_2_0_47), .A2(n_2_0_16), .ZN(n_2_404));
   NOR2_X1 i_2_0_576 (.A1(n_2_0_47), .A2(n_2_0_17), .ZN(n_2_405));
   NOR2_X1 i_2_0_577 (.A1(n_2_0_47), .A2(n_2_0_18), .ZN(n_2_406));
   NOR2_X1 i_2_0_578 (.A1(n_2_0_47), .A2(n_2_0_19), .ZN(n_2_407));
   NOR2_X1 i_2_0_579 (.A1(n_2_0_47), .A2(n_2_0_20), .ZN(n_2_408));
   NOR2_X1 i_2_0_580 (.A1(n_2_0_47), .A2(n_2_0_21), .ZN(n_2_409));
   NOR2_X1 i_2_0_581 (.A1(n_2_0_47), .A2(n_2_0_22), .ZN(n_2_410));
   NOR2_X1 i_2_0_582 (.A1(n_2_0_47), .A2(n_2_0_23), .ZN(n_2_411));
   NOR2_X1 i_2_0_583 (.A1(n_2_0_47), .A2(n_2_0_24), .ZN(n_2_412));
   NOR2_X1 i_2_0_584 (.A1(n_2_0_47), .A2(n_2_0_25), .ZN(n_2_413));
   NOR2_X1 i_2_0_585 (.A1(n_2_0_47), .A2(n_2_0_26), .ZN(n_2_414));
   NOR2_X1 i_2_0_586 (.A1(n_2_0_47), .A2(n_2_0_27), .ZN(n_2_415));
   NOR2_X1 i_2_0_587 (.A1(n_2_0_47), .A2(n_2_0_28), .ZN(n_2_416));
   NOR2_X1 i_2_0_588 (.A1(n_2_0_47), .A2(n_2_0_29), .ZN(n_2_417));
   NOR2_X1 i_2_0_589 (.A1(n_2_0_47), .A2(n_2_0_30), .ZN(n_2_418));
   NOR2_X1 i_2_0_590 (.A1(n_2_0_47), .A2(n_2_0_31), .ZN(n_2_419));
   NOR2_X1 i_2_0_591 (.A1(n_2_0_47), .A2(n_2_0_32), .ZN(n_2_420));
   INV_X1 i_2_0_592 (.A(n_802), .ZN(n_2_0_48));
   NOR2_X1 i_2_0_593 (.A1(n_2_0_48), .A2(n_2_0_1), .ZN(n_2_421));
   NOR2_X1 i_2_0_594 (.A1(n_2_0_48), .A2(n_2_0_2), .ZN(n_2_422));
   NOR2_X1 i_2_0_595 (.A1(n_2_0_48), .A2(n_2_0_3), .ZN(n_2_423));
   NOR2_X1 i_2_0_596 (.A1(n_2_0_48), .A2(n_2_0_4), .ZN(n_2_424));
   NOR2_X1 i_2_0_597 (.A1(n_2_0_48), .A2(n_2_0_5), .ZN(n_2_425));
   NOR2_X1 i_2_0_598 (.A1(n_2_0_48), .A2(n_2_0_6), .ZN(n_2_426));
   NOR2_X1 i_2_0_599 (.A1(n_2_0_48), .A2(n_2_0_7), .ZN(n_2_427));
   NOR2_X1 i_2_0_600 (.A1(n_2_0_48), .A2(n_2_0_8), .ZN(n_2_428));
   NOR2_X1 i_2_0_601 (.A1(n_2_0_48), .A2(n_2_0_9), .ZN(n_2_429));
   NOR2_X1 i_2_0_602 (.A1(n_2_0_48), .A2(n_2_0_10), .ZN(n_2_430));
   NOR2_X1 i_2_0_603 (.A1(n_2_0_48), .A2(n_2_0_11), .ZN(n_2_431));
   NOR2_X1 i_2_0_604 (.A1(n_2_0_48), .A2(n_2_0_12), .ZN(n_2_432));
   NOR2_X1 i_2_0_605 (.A1(n_2_0_48), .A2(n_2_0_13), .ZN(n_2_433));
   NOR2_X1 i_2_0_606 (.A1(n_2_0_48), .A2(n_2_0_14), .ZN(n_2_434));
   NOR2_X1 i_2_0_607 (.A1(n_2_0_48), .A2(n_2_0_15), .ZN(n_2_435));
   NOR2_X1 i_2_0_608 (.A1(n_2_0_48), .A2(n_2_0_16), .ZN(n_2_436));
   NOR2_X1 i_2_0_609 (.A1(n_2_0_48), .A2(n_2_0_17), .ZN(n_2_437));
   NOR2_X1 i_2_0_610 (.A1(n_2_0_48), .A2(n_2_0_18), .ZN(n_2_438));
   NOR2_X1 i_2_0_611 (.A1(n_2_0_48), .A2(n_2_0_19), .ZN(n_2_439));
   NOR2_X1 i_2_0_612 (.A1(n_2_0_48), .A2(n_2_0_20), .ZN(n_2_440));
   NOR2_X1 i_2_0_613 (.A1(n_2_0_48), .A2(n_2_0_21), .ZN(n_2_441));
   NOR2_X1 i_2_0_614 (.A1(n_2_0_48), .A2(n_2_0_22), .ZN(n_2_442));
   NOR2_X1 i_2_0_615 (.A1(n_2_0_48), .A2(n_2_0_23), .ZN(n_2_443));
   NOR2_X1 i_2_0_616 (.A1(n_2_0_48), .A2(n_2_0_24), .ZN(n_2_444));
   NOR2_X1 i_2_0_617 (.A1(n_2_0_48), .A2(n_2_0_25), .ZN(n_2_445));
   NOR2_X1 i_2_0_618 (.A1(n_2_0_48), .A2(n_2_0_26), .ZN(n_2_446));
   NOR2_X1 i_2_0_619 (.A1(n_2_0_48), .A2(n_2_0_27), .ZN(n_2_447));
   NOR2_X1 i_2_0_620 (.A1(n_2_0_48), .A2(n_2_0_28), .ZN(n_2_448));
   NOR2_X1 i_2_0_621 (.A1(n_2_0_48), .A2(n_2_0_29), .ZN(n_2_449));
   NOR2_X1 i_2_0_622 (.A1(n_2_0_48), .A2(n_2_0_30), .ZN(n_2_450));
   NOR2_X1 i_2_0_623 (.A1(n_2_0_48), .A2(n_2_0_31), .ZN(n_2_451));
   NOR2_X1 i_2_0_624 (.A1(n_2_0_48), .A2(n_2_0_32), .ZN(n_2_452));
   INV_X1 i_2_0_625 (.A(n_801), .ZN(n_2_0_49));
   NOR2_X1 i_2_0_626 (.A1(n_2_0_49), .A2(n_2_0_1), .ZN(n_2_453));
   NOR2_X1 i_2_0_627 (.A1(n_2_0_49), .A2(n_2_0_2), .ZN(n_2_454));
   NOR2_X1 i_2_0_628 (.A1(n_2_0_49), .A2(n_2_0_3), .ZN(n_2_455));
   NOR2_X1 i_2_0_629 (.A1(n_2_0_49), .A2(n_2_0_4), .ZN(n_2_456));
   NOR2_X1 i_2_0_630 (.A1(n_2_0_49), .A2(n_2_0_5), .ZN(n_2_457));
   NOR2_X1 i_2_0_631 (.A1(n_2_0_49), .A2(n_2_0_6), .ZN(n_2_458));
   NOR2_X1 i_2_0_632 (.A1(n_2_0_49), .A2(n_2_0_7), .ZN(n_2_459));
   NOR2_X1 i_2_0_633 (.A1(n_2_0_49), .A2(n_2_0_8), .ZN(n_2_460));
   NOR2_X1 i_2_0_634 (.A1(n_2_0_49), .A2(n_2_0_9), .ZN(n_2_461));
   NOR2_X1 i_2_0_635 (.A1(n_2_0_49), .A2(n_2_0_10), .ZN(n_2_462));
   NOR2_X1 i_2_0_636 (.A1(n_2_0_49), .A2(n_2_0_11), .ZN(n_2_463));
   NOR2_X1 i_2_0_637 (.A1(n_2_0_49), .A2(n_2_0_12), .ZN(n_2_464));
   NOR2_X1 i_2_0_638 (.A1(n_2_0_49), .A2(n_2_0_13), .ZN(n_2_465));
   NOR2_X1 i_2_0_639 (.A1(n_2_0_49), .A2(n_2_0_14), .ZN(n_2_466));
   NOR2_X1 i_2_0_640 (.A1(n_2_0_49), .A2(n_2_0_15), .ZN(n_2_467));
   NOR2_X1 i_2_0_641 (.A1(n_2_0_49), .A2(n_2_0_16), .ZN(n_2_468));
   NOR2_X1 i_2_0_642 (.A1(n_2_0_49), .A2(n_2_0_17), .ZN(n_2_469));
   NOR2_X1 i_2_0_643 (.A1(n_2_0_49), .A2(n_2_0_18), .ZN(n_2_470));
   NOR2_X1 i_2_0_644 (.A1(n_2_0_49), .A2(n_2_0_19), .ZN(n_2_471));
   NOR2_X1 i_2_0_645 (.A1(n_2_0_49), .A2(n_2_0_20), .ZN(n_2_472));
   NOR2_X1 i_2_0_646 (.A1(n_2_0_49), .A2(n_2_0_21), .ZN(n_2_473));
   NOR2_X1 i_2_0_647 (.A1(n_2_0_49), .A2(n_2_0_22), .ZN(n_2_474));
   NOR2_X1 i_2_0_648 (.A1(n_2_0_49), .A2(n_2_0_23), .ZN(n_2_475));
   NOR2_X1 i_2_0_649 (.A1(n_2_0_49), .A2(n_2_0_24), .ZN(n_2_476));
   NOR2_X1 i_2_0_650 (.A1(n_2_0_49), .A2(n_2_0_25), .ZN(n_2_477));
   NOR2_X1 i_2_0_651 (.A1(n_2_0_49), .A2(n_2_0_26), .ZN(n_2_478));
   NOR2_X1 i_2_0_652 (.A1(n_2_0_49), .A2(n_2_0_27), .ZN(n_2_479));
   NOR2_X1 i_2_0_653 (.A1(n_2_0_49), .A2(n_2_0_28), .ZN(n_2_480));
   NOR2_X1 i_2_0_654 (.A1(n_2_0_49), .A2(n_2_0_29), .ZN(n_2_481));
   NOR2_X1 i_2_0_655 (.A1(n_2_0_49), .A2(n_2_0_30), .ZN(n_2_482));
   NOR2_X1 i_2_0_656 (.A1(n_2_0_49), .A2(n_2_0_31), .ZN(n_2_483));
   NOR2_X1 i_2_0_657 (.A1(n_2_0_49), .A2(n_2_0_32), .ZN(n_2_484));
   INV_X1 i_2_0_658 (.A(n_800), .ZN(n_2_0_50));
   NOR2_X1 i_2_0_659 (.A1(n_2_0_50), .A2(n_2_0_1), .ZN(n_2_485));
   NOR2_X1 i_2_0_660 (.A1(n_2_0_50), .A2(n_2_0_2), .ZN(n_2_486));
   NOR2_X1 i_2_0_661 (.A1(n_2_0_50), .A2(n_2_0_3), .ZN(n_2_487));
   NOR2_X1 i_2_0_662 (.A1(n_2_0_50), .A2(n_2_0_4), .ZN(n_2_488));
   NOR2_X1 i_2_0_663 (.A1(n_2_0_50), .A2(n_2_0_5), .ZN(n_2_489));
   NOR2_X1 i_2_0_664 (.A1(n_2_0_50), .A2(n_2_0_6), .ZN(n_2_490));
   NOR2_X1 i_2_0_665 (.A1(n_2_0_50), .A2(n_2_0_7), .ZN(n_2_491));
   NOR2_X1 i_2_0_666 (.A1(n_2_0_50), .A2(n_2_0_8), .ZN(n_2_492));
   NOR2_X1 i_2_0_667 (.A1(n_2_0_50), .A2(n_2_0_9), .ZN(n_2_493));
   NOR2_X1 i_2_0_668 (.A1(n_2_0_50), .A2(n_2_0_10), .ZN(n_2_494));
   NOR2_X1 i_2_0_669 (.A1(n_2_0_50), .A2(n_2_0_11), .ZN(n_2_495));
   NOR2_X1 i_2_0_670 (.A1(n_2_0_50), .A2(n_2_0_12), .ZN(n_2_496));
   NOR2_X1 i_2_0_671 (.A1(n_2_0_50), .A2(n_2_0_13), .ZN(n_2_497));
   NOR2_X1 i_2_0_672 (.A1(n_2_0_50), .A2(n_2_0_14), .ZN(n_2_498));
   NOR2_X1 i_2_0_673 (.A1(n_2_0_50), .A2(n_2_0_15), .ZN(n_2_499));
   NOR2_X1 i_2_0_674 (.A1(n_2_0_50), .A2(n_2_0_16), .ZN(n_2_500));
   NOR2_X1 i_2_0_675 (.A1(n_2_0_50), .A2(n_2_0_17), .ZN(n_2_501));
   NOR2_X1 i_2_0_676 (.A1(n_2_0_50), .A2(n_2_0_18), .ZN(n_2_502));
   NOR2_X1 i_2_0_677 (.A1(n_2_0_50), .A2(n_2_0_19), .ZN(n_2_503));
   NOR2_X1 i_2_0_678 (.A1(n_2_0_50), .A2(n_2_0_20), .ZN(n_2_504));
   NOR2_X1 i_2_0_679 (.A1(n_2_0_50), .A2(n_2_0_21), .ZN(n_2_505));
   NOR2_X1 i_2_0_680 (.A1(n_2_0_50), .A2(n_2_0_22), .ZN(n_2_506));
   NOR2_X1 i_2_0_681 (.A1(n_2_0_50), .A2(n_2_0_23), .ZN(n_2_507));
   NOR2_X1 i_2_0_682 (.A1(n_2_0_50), .A2(n_2_0_24), .ZN(n_2_508));
   NOR2_X1 i_2_0_683 (.A1(n_2_0_50), .A2(n_2_0_25), .ZN(n_2_509));
   NOR2_X1 i_2_0_684 (.A1(n_2_0_50), .A2(n_2_0_26), .ZN(n_2_510));
   NOR2_X1 i_2_0_685 (.A1(n_2_0_50), .A2(n_2_0_27), .ZN(n_2_511));
   NOR2_X1 i_2_0_686 (.A1(n_2_0_50), .A2(n_2_0_28), .ZN(n_2_512));
   NOR2_X1 i_2_0_687 (.A1(n_2_0_50), .A2(n_2_0_29), .ZN(n_2_513));
   NOR2_X1 i_2_0_688 (.A1(n_2_0_50), .A2(n_2_0_30), .ZN(n_2_514));
   NOR2_X1 i_2_0_689 (.A1(n_2_0_50), .A2(n_2_0_31), .ZN(n_2_515));
   NOR2_X1 i_2_0_690 (.A1(n_2_0_50), .A2(n_2_0_32), .ZN(n_2_516));
   INV_X1 i_2_0_691 (.A(n_799), .ZN(n_2_0_51));
   NOR2_X1 i_2_0_692 (.A1(n_2_0_51), .A2(n_2_0_1), .ZN(n_2_517));
   NOR2_X1 i_2_0_693 (.A1(n_2_0_51), .A2(n_2_0_2), .ZN(n_2_518));
   NOR2_X1 i_2_0_694 (.A1(n_2_0_51), .A2(n_2_0_3), .ZN(n_2_519));
   NOR2_X1 i_2_0_695 (.A1(n_2_0_51), .A2(n_2_0_4), .ZN(n_2_520));
   NOR2_X1 i_2_0_696 (.A1(n_2_0_51), .A2(n_2_0_5), .ZN(n_2_521));
   NOR2_X1 i_2_0_697 (.A1(n_2_0_51), .A2(n_2_0_6), .ZN(n_2_522));
   NOR2_X1 i_2_0_698 (.A1(n_2_0_51), .A2(n_2_0_7), .ZN(n_2_523));
   NOR2_X1 i_2_0_699 (.A1(n_2_0_51), .A2(n_2_0_8), .ZN(n_2_524));
   NOR2_X1 i_2_0_700 (.A1(n_2_0_51), .A2(n_2_0_9), .ZN(n_2_525));
   NOR2_X1 i_2_0_701 (.A1(n_2_0_51), .A2(n_2_0_10), .ZN(n_2_526));
   NOR2_X1 i_2_0_702 (.A1(n_2_0_51), .A2(n_2_0_11), .ZN(n_2_527));
   NOR2_X1 i_2_0_703 (.A1(n_2_0_51), .A2(n_2_0_12), .ZN(n_2_528));
   NOR2_X1 i_2_0_704 (.A1(n_2_0_51), .A2(n_2_0_13), .ZN(n_2_529));
   NOR2_X1 i_2_0_705 (.A1(n_2_0_51), .A2(n_2_0_14), .ZN(n_2_530));
   NOR2_X1 i_2_0_706 (.A1(n_2_0_51), .A2(n_2_0_15), .ZN(n_2_531));
   NOR2_X1 i_2_0_707 (.A1(n_2_0_51), .A2(n_2_0_16), .ZN(n_2_532));
   NOR2_X1 i_2_0_708 (.A1(n_2_0_51), .A2(n_2_0_17), .ZN(n_2_533));
   NOR2_X1 i_2_0_709 (.A1(n_2_0_51), .A2(n_2_0_18), .ZN(n_2_534));
   NOR2_X1 i_2_0_710 (.A1(n_2_0_51), .A2(n_2_0_19), .ZN(n_2_535));
   NOR2_X1 i_2_0_711 (.A1(n_2_0_51), .A2(n_2_0_20), .ZN(n_2_536));
   NOR2_X1 i_2_0_712 (.A1(n_2_0_51), .A2(n_2_0_21), .ZN(n_2_537));
   NOR2_X1 i_2_0_713 (.A1(n_2_0_51), .A2(n_2_0_22), .ZN(n_2_538));
   NOR2_X1 i_2_0_714 (.A1(n_2_0_51), .A2(n_2_0_23), .ZN(n_2_539));
   NOR2_X1 i_2_0_715 (.A1(n_2_0_51), .A2(n_2_0_24), .ZN(n_2_540));
   NOR2_X1 i_2_0_716 (.A1(n_2_0_51), .A2(n_2_0_25), .ZN(n_2_541));
   NOR2_X1 i_2_0_717 (.A1(n_2_0_51), .A2(n_2_0_26), .ZN(n_2_542));
   NOR2_X1 i_2_0_718 (.A1(n_2_0_51), .A2(n_2_0_27), .ZN(n_2_543));
   NOR2_X1 i_2_0_719 (.A1(n_2_0_51), .A2(n_2_0_28), .ZN(n_2_544));
   NOR2_X1 i_2_0_720 (.A1(n_2_0_51), .A2(n_2_0_29), .ZN(n_2_545));
   NOR2_X1 i_2_0_721 (.A1(n_2_0_51), .A2(n_2_0_30), .ZN(n_2_546));
   NOR2_X1 i_2_0_722 (.A1(n_2_0_51), .A2(n_2_0_31), .ZN(n_2_547));
   NOR2_X1 i_2_0_723 (.A1(n_2_0_51), .A2(n_2_0_32), .ZN(n_2_548));
   INV_X1 i_2_0_724 (.A(n_798), .ZN(n_2_0_52));
   NOR2_X1 i_2_0_725 (.A1(n_2_0_52), .A2(n_2_0_1), .ZN(n_2_549));
   NOR2_X1 i_2_0_726 (.A1(n_2_0_52), .A2(n_2_0_2), .ZN(n_2_550));
   NOR2_X1 i_2_0_727 (.A1(n_2_0_52), .A2(n_2_0_3), .ZN(n_2_551));
   NOR2_X1 i_2_0_728 (.A1(n_2_0_52), .A2(n_2_0_4), .ZN(n_2_552));
   NOR2_X1 i_2_0_729 (.A1(n_2_0_52), .A2(n_2_0_5), .ZN(n_2_553));
   NOR2_X1 i_2_0_730 (.A1(n_2_0_52), .A2(n_2_0_6), .ZN(n_2_554));
   NOR2_X1 i_2_0_731 (.A1(n_2_0_52), .A2(n_2_0_7), .ZN(n_2_555));
   NOR2_X1 i_2_0_732 (.A1(n_2_0_52), .A2(n_2_0_8), .ZN(n_2_556));
   NOR2_X1 i_2_0_733 (.A1(n_2_0_52), .A2(n_2_0_9), .ZN(n_2_557));
   NOR2_X1 i_2_0_734 (.A1(n_2_0_52), .A2(n_2_0_10), .ZN(n_2_558));
   NOR2_X1 i_2_0_735 (.A1(n_2_0_52), .A2(n_2_0_11), .ZN(n_2_559));
   NOR2_X1 i_2_0_736 (.A1(n_2_0_52), .A2(n_2_0_12), .ZN(n_2_560));
   NOR2_X1 i_2_0_737 (.A1(n_2_0_52), .A2(n_2_0_13), .ZN(n_2_561));
   NOR2_X1 i_2_0_738 (.A1(n_2_0_52), .A2(n_2_0_14), .ZN(n_2_562));
   NOR2_X1 i_2_0_739 (.A1(n_2_0_52), .A2(n_2_0_15), .ZN(n_2_563));
   NOR2_X1 i_2_0_740 (.A1(n_2_0_52), .A2(n_2_0_16), .ZN(n_2_564));
   NOR2_X1 i_2_0_741 (.A1(n_2_0_52), .A2(n_2_0_17), .ZN(n_2_565));
   NOR2_X1 i_2_0_742 (.A1(n_2_0_52), .A2(n_2_0_18), .ZN(n_2_566));
   NOR2_X1 i_2_0_743 (.A1(n_2_0_52), .A2(n_2_0_19), .ZN(n_2_567));
   NOR2_X1 i_2_0_744 (.A1(n_2_0_52), .A2(n_2_0_20), .ZN(n_2_568));
   NOR2_X1 i_2_0_745 (.A1(n_2_0_52), .A2(n_2_0_21), .ZN(n_2_569));
   NOR2_X1 i_2_0_746 (.A1(n_2_0_52), .A2(n_2_0_22), .ZN(n_2_570));
   NOR2_X1 i_2_0_747 (.A1(n_2_0_52), .A2(n_2_0_23), .ZN(n_2_571));
   NOR2_X1 i_2_0_748 (.A1(n_2_0_52), .A2(n_2_0_24), .ZN(n_2_572));
   NOR2_X1 i_2_0_749 (.A1(n_2_0_52), .A2(n_2_0_25), .ZN(n_2_573));
   NOR2_X1 i_2_0_750 (.A1(n_2_0_52), .A2(n_2_0_26), .ZN(n_2_574));
   NOR2_X1 i_2_0_751 (.A1(n_2_0_52), .A2(n_2_0_27), .ZN(n_2_575));
   NOR2_X1 i_2_0_752 (.A1(n_2_0_52), .A2(n_2_0_28), .ZN(n_2_576));
   NOR2_X1 i_2_0_753 (.A1(n_2_0_52), .A2(n_2_0_29), .ZN(n_2_577));
   NOR2_X1 i_2_0_754 (.A1(n_2_0_52), .A2(n_2_0_30), .ZN(n_2_578));
   NOR2_X1 i_2_0_755 (.A1(n_2_0_52), .A2(n_2_0_31), .ZN(n_2_579));
   NOR2_X1 i_2_0_756 (.A1(n_2_0_52), .A2(n_2_0_32), .ZN(n_2_580));
   INV_X1 i_2_0_757 (.A(n_797), .ZN(n_2_0_53));
   NOR2_X1 i_2_0_758 (.A1(n_2_0_53), .A2(n_2_0_1), .ZN(n_2_581));
   NOR2_X1 i_2_0_759 (.A1(n_2_0_53), .A2(n_2_0_2), .ZN(n_2_582));
   NOR2_X1 i_2_0_760 (.A1(n_2_0_53), .A2(n_2_0_3), .ZN(n_2_583));
   NOR2_X1 i_2_0_761 (.A1(n_2_0_53), .A2(n_2_0_4), .ZN(n_2_584));
   NOR2_X1 i_2_0_762 (.A1(n_2_0_53), .A2(n_2_0_5), .ZN(n_2_585));
   NOR2_X1 i_2_0_763 (.A1(n_2_0_53), .A2(n_2_0_6), .ZN(n_2_586));
   NOR2_X1 i_2_0_764 (.A1(n_2_0_53), .A2(n_2_0_7), .ZN(n_2_587));
   NOR2_X1 i_2_0_765 (.A1(n_2_0_53), .A2(n_2_0_8), .ZN(n_2_588));
   NOR2_X1 i_2_0_766 (.A1(n_2_0_53), .A2(n_2_0_9), .ZN(n_2_589));
   NOR2_X1 i_2_0_767 (.A1(n_2_0_53), .A2(n_2_0_10), .ZN(n_2_590));
   NOR2_X1 i_2_0_768 (.A1(n_2_0_53), .A2(n_2_0_11), .ZN(n_2_591));
   NOR2_X1 i_2_0_769 (.A1(n_2_0_53), .A2(n_2_0_12), .ZN(n_2_592));
   NOR2_X1 i_2_0_770 (.A1(n_2_0_53), .A2(n_2_0_13), .ZN(n_2_593));
   NOR2_X1 i_2_0_771 (.A1(n_2_0_53), .A2(n_2_0_14), .ZN(n_2_594));
   NOR2_X1 i_2_0_772 (.A1(n_2_0_53), .A2(n_2_0_15), .ZN(n_2_595));
   NOR2_X1 i_2_0_773 (.A1(n_2_0_53), .A2(n_2_0_16), .ZN(n_2_596));
   NOR2_X1 i_2_0_774 (.A1(n_2_0_53), .A2(n_2_0_17), .ZN(n_2_597));
   NOR2_X1 i_2_0_775 (.A1(n_2_0_53), .A2(n_2_0_18), .ZN(n_2_598));
   NOR2_X1 i_2_0_776 (.A1(n_2_0_53), .A2(n_2_0_19), .ZN(n_2_599));
   NOR2_X1 i_2_0_777 (.A1(n_2_0_53), .A2(n_2_0_20), .ZN(n_2_600));
   NOR2_X1 i_2_0_778 (.A1(n_2_0_53), .A2(n_2_0_21), .ZN(n_2_601));
   NOR2_X1 i_2_0_779 (.A1(n_2_0_53), .A2(n_2_0_22), .ZN(n_2_602));
   NOR2_X1 i_2_0_780 (.A1(n_2_0_53), .A2(n_2_0_23), .ZN(n_2_603));
   NOR2_X1 i_2_0_781 (.A1(n_2_0_53), .A2(n_2_0_24), .ZN(n_2_604));
   NOR2_X1 i_2_0_782 (.A1(n_2_0_53), .A2(n_2_0_25), .ZN(n_2_605));
   NOR2_X1 i_2_0_783 (.A1(n_2_0_53), .A2(n_2_0_26), .ZN(n_2_606));
   NOR2_X1 i_2_0_784 (.A1(n_2_0_53), .A2(n_2_0_27), .ZN(n_2_607));
   NOR2_X1 i_2_0_785 (.A1(n_2_0_53), .A2(n_2_0_28), .ZN(n_2_608));
   NOR2_X1 i_2_0_786 (.A1(n_2_0_53), .A2(n_2_0_29), .ZN(n_2_609));
   NOR2_X1 i_2_0_787 (.A1(n_2_0_53), .A2(n_2_0_30), .ZN(n_2_610));
   NOR2_X1 i_2_0_788 (.A1(n_2_0_53), .A2(n_2_0_31), .ZN(n_2_611));
   NOR2_X1 i_2_0_789 (.A1(n_2_0_53), .A2(n_2_0_32), .ZN(n_2_612));
   INV_X1 i_2_0_790 (.A(n_796), .ZN(n_2_0_54));
   NOR2_X1 i_2_0_791 (.A1(n_2_0_54), .A2(n_2_0_1), .ZN(n_164));
   NOR2_X1 i_2_0_792 (.A1(n_2_0_54), .A2(n_2_0_2), .ZN(n_2_613));
   NOR2_X1 i_2_0_793 (.A1(n_2_0_54), .A2(n_2_0_3), .ZN(n_2_614));
   NOR2_X1 i_2_0_794 (.A1(n_2_0_54), .A2(n_2_0_4), .ZN(n_2_615));
   NOR2_X1 i_2_0_795 (.A1(n_2_0_54), .A2(n_2_0_5), .ZN(n_2_616));
   NOR2_X1 i_2_0_796 (.A1(n_2_0_54), .A2(n_2_0_6), .ZN(n_2_617));
   NOR2_X1 i_2_0_797 (.A1(n_2_0_54), .A2(n_2_0_7), .ZN(n_2_618));
   NOR2_X1 i_2_0_798 (.A1(n_2_0_54), .A2(n_2_0_8), .ZN(n_2_619));
   NOR2_X1 i_2_0_799 (.A1(n_2_0_54), .A2(n_2_0_9), .ZN(n_2_620));
   NOR2_X1 i_2_0_800 (.A1(n_2_0_54), .A2(n_2_0_10), .ZN(n_2_621));
   NOR2_X1 i_2_0_801 (.A1(n_2_0_54), .A2(n_2_0_11), .ZN(n_2_622));
   NOR2_X1 i_2_0_802 (.A1(n_2_0_54), .A2(n_2_0_12), .ZN(n_2_623));
   NOR2_X1 i_2_0_803 (.A1(n_2_0_54), .A2(n_2_0_13), .ZN(n_2_624));
   NOR2_X1 i_2_0_804 (.A1(n_2_0_54), .A2(n_2_0_14), .ZN(n_2_625));
   NOR2_X1 i_2_0_805 (.A1(n_2_0_54), .A2(n_2_0_15), .ZN(n_2_626));
   NOR2_X1 i_2_0_806 (.A1(n_2_0_54), .A2(n_2_0_16), .ZN(n_2_627));
   NOR2_X1 i_2_0_807 (.A1(n_2_0_54), .A2(n_2_0_17), .ZN(n_2_628));
   NOR2_X1 i_2_0_808 (.A1(n_2_0_54), .A2(n_2_0_18), .ZN(n_2_629));
   NOR2_X1 i_2_0_809 (.A1(n_2_0_54), .A2(n_2_0_19), .ZN(n_2_630));
   NOR2_X1 i_2_0_810 (.A1(n_2_0_54), .A2(n_2_0_20), .ZN(n_2_631));
   NOR2_X1 i_2_0_811 (.A1(n_2_0_54), .A2(n_2_0_21), .ZN(n_2_632));
   NOR2_X1 i_2_0_812 (.A1(n_2_0_54), .A2(n_2_0_22), .ZN(n_2_633));
   NOR2_X1 i_2_0_813 (.A1(n_2_0_54), .A2(n_2_0_23), .ZN(n_2_634));
   NOR2_X1 i_2_0_814 (.A1(n_2_0_54), .A2(n_2_0_24), .ZN(n_2_635));
   NOR2_X1 i_2_0_815 (.A1(n_2_0_54), .A2(n_2_0_25), .ZN(n_2_636));
   NOR2_X1 i_2_0_816 (.A1(n_2_0_54), .A2(n_2_0_26), .ZN(n_2_637));
   NOR2_X1 i_2_0_817 (.A1(n_2_0_54), .A2(n_2_0_27), .ZN(n_2_638));
   NOR2_X1 i_2_0_818 (.A1(n_2_0_54), .A2(n_2_0_28), .ZN(n_2_639));
   NOR2_X1 i_2_0_819 (.A1(n_2_0_54), .A2(n_2_0_29), .ZN(n_2_640));
   NOR2_X1 i_2_0_820 (.A1(n_2_0_54), .A2(n_2_0_30), .ZN(n_2_641));
   NOR2_X1 i_2_0_821 (.A1(n_2_0_54), .A2(n_2_0_31), .ZN(n_2_642));
   NOR2_X1 i_2_0_822 (.A1(n_2_0_54), .A2(n_2_0_32), .ZN(n_2_643));
   INV_X1 i_2_0_823 (.A(n_795), .ZN(n_2_0_55));
   NOR2_X1 i_2_0_824 (.A1(n_2_0_55), .A2(n_2_0_1), .ZN(n_2_644));
   NOR2_X1 i_2_0_825 (.A1(n_2_0_55), .A2(n_2_0_2), .ZN(n_2_645));
   NOR2_X1 i_2_0_826 (.A1(n_2_0_55), .A2(n_2_0_3), .ZN(n_2_646));
   NOR2_X1 i_2_0_827 (.A1(n_2_0_55), .A2(n_2_0_4), .ZN(n_2_647));
   NOR2_X1 i_2_0_828 (.A1(n_2_0_55), .A2(n_2_0_5), .ZN(n_2_648));
   NOR2_X1 i_2_0_829 (.A1(n_2_0_55), .A2(n_2_0_6), .ZN(n_2_649));
   NOR2_X1 i_2_0_830 (.A1(n_2_0_55), .A2(n_2_0_7), .ZN(n_2_650));
   NOR2_X1 i_2_0_831 (.A1(n_2_0_55), .A2(n_2_0_8), .ZN(n_2_651));
   NOR2_X1 i_2_0_832 (.A1(n_2_0_55), .A2(n_2_0_9), .ZN(n_2_652));
   NOR2_X1 i_2_0_833 (.A1(n_2_0_55), .A2(n_2_0_10), .ZN(n_2_653));
   NOR2_X1 i_2_0_834 (.A1(n_2_0_55), .A2(n_2_0_11), .ZN(n_2_654));
   NOR2_X1 i_2_0_835 (.A1(n_2_0_55), .A2(n_2_0_12), .ZN(n_2_655));
   NOR2_X1 i_2_0_836 (.A1(n_2_0_55), .A2(n_2_0_13), .ZN(n_2_656));
   NOR2_X1 i_2_0_837 (.A1(n_2_0_55), .A2(n_2_0_14), .ZN(n_2_657));
   NOR2_X1 i_2_0_838 (.A1(n_2_0_55), .A2(n_2_0_15), .ZN(n_2_658));
   NOR2_X1 i_2_0_839 (.A1(n_2_0_55), .A2(n_2_0_16), .ZN(n_2_659));
   NOR2_X1 i_2_0_840 (.A1(n_2_0_55), .A2(n_2_0_17), .ZN(n_2_660));
   NOR2_X1 i_2_0_841 (.A1(n_2_0_55), .A2(n_2_0_18), .ZN(n_2_661));
   NOR2_X1 i_2_0_842 (.A1(n_2_0_55), .A2(n_2_0_19), .ZN(n_2_662));
   NOR2_X1 i_2_0_843 (.A1(n_2_0_55), .A2(n_2_0_20), .ZN(n_2_663));
   NOR2_X1 i_2_0_844 (.A1(n_2_0_55), .A2(n_2_0_21), .ZN(n_2_664));
   NOR2_X1 i_2_0_845 (.A1(n_2_0_55), .A2(n_2_0_22), .ZN(n_2_665));
   NOR2_X1 i_2_0_846 (.A1(n_2_0_55), .A2(n_2_0_23), .ZN(n_2_666));
   NOR2_X1 i_2_0_847 (.A1(n_2_0_55), .A2(n_2_0_24), .ZN(n_2_667));
   NOR2_X1 i_2_0_848 (.A1(n_2_0_55), .A2(n_2_0_25), .ZN(n_2_668));
   NOR2_X1 i_2_0_849 (.A1(n_2_0_55), .A2(n_2_0_26), .ZN(n_2_669));
   NOR2_X1 i_2_0_850 (.A1(n_2_0_55), .A2(n_2_0_27), .ZN(n_2_670));
   NOR2_X1 i_2_0_851 (.A1(n_2_0_55), .A2(n_2_0_28), .ZN(n_2_671));
   NOR2_X1 i_2_0_852 (.A1(n_2_0_55), .A2(n_2_0_29), .ZN(n_2_672));
   NOR2_X1 i_2_0_853 (.A1(n_2_0_55), .A2(n_2_0_30), .ZN(n_2_673));
   NOR2_X1 i_2_0_854 (.A1(n_2_0_55), .A2(n_2_0_31), .ZN(n_2_674));
   NOR2_X1 i_2_0_855 (.A1(n_2_0_55), .A2(n_2_0_32), .ZN(n_2_675));
   INV_X1 i_2_0_856 (.A(n_794), .ZN(n_2_0_56));
   NOR2_X1 i_2_0_857 (.A1(n_2_0_56), .A2(n_2_0_1), .ZN(n_2_676));
   NOR2_X1 i_2_0_858 (.A1(n_2_0_56), .A2(n_2_0_2), .ZN(n_2_677));
   NOR2_X1 i_2_0_859 (.A1(n_2_0_56), .A2(n_2_0_3), .ZN(n_2_678));
   NOR2_X1 i_2_0_860 (.A1(n_2_0_56), .A2(n_2_0_4), .ZN(n_2_679));
   NOR2_X1 i_2_0_861 (.A1(n_2_0_56), .A2(n_2_0_5), .ZN(n_2_680));
   NOR2_X1 i_2_0_862 (.A1(n_2_0_56), .A2(n_2_0_6), .ZN(n_2_681));
   NOR2_X1 i_2_0_863 (.A1(n_2_0_56), .A2(n_2_0_7), .ZN(n_2_682));
   NOR2_X1 i_2_0_864 (.A1(n_2_0_56), .A2(n_2_0_8), .ZN(n_2_683));
   NOR2_X1 i_2_0_865 (.A1(n_2_0_56), .A2(n_2_0_9), .ZN(n_2_684));
   NOR2_X1 i_2_0_866 (.A1(n_2_0_56), .A2(n_2_0_10), .ZN(n_2_685));
   NOR2_X1 i_2_0_867 (.A1(n_2_0_56), .A2(n_2_0_11), .ZN(n_2_686));
   NOR2_X1 i_2_0_868 (.A1(n_2_0_56), .A2(n_2_0_12), .ZN(n_2_687));
   NOR2_X1 i_2_0_869 (.A1(n_2_0_56), .A2(n_2_0_13), .ZN(n_2_688));
   NOR2_X1 i_2_0_870 (.A1(n_2_0_56), .A2(n_2_0_14), .ZN(n_2_689));
   NOR2_X1 i_2_0_871 (.A1(n_2_0_56), .A2(n_2_0_15), .ZN(n_2_690));
   NOR2_X1 i_2_0_872 (.A1(n_2_0_56), .A2(n_2_0_16), .ZN(n_2_691));
   NOR2_X1 i_2_0_873 (.A1(n_2_0_56), .A2(n_2_0_17), .ZN(n_2_692));
   NOR2_X1 i_2_0_874 (.A1(n_2_0_56), .A2(n_2_0_18), .ZN(n_2_693));
   NOR2_X1 i_2_0_875 (.A1(n_2_0_56), .A2(n_2_0_19), .ZN(n_2_694));
   NOR2_X1 i_2_0_876 (.A1(n_2_0_56), .A2(n_2_0_20), .ZN(n_2_695));
   NOR2_X1 i_2_0_877 (.A1(n_2_0_56), .A2(n_2_0_21), .ZN(n_2_696));
   NOR2_X1 i_2_0_878 (.A1(n_2_0_56), .A2(n_2_0_22), .ZN(n_2_697));
   NOR2_X1 i_2_0_879 (.A1(n_2_0_56), .A2(n_2_0_23), .ZN(n_2_698));
   NOR2_X1 i_2_0_880 (.A1(n_2_0_56), .A2(n_2_0_24), .ZN(n_2_699));
   NOR2_X1 i_2_0_881 (.A1(n_2_0_56), .A2(n_2_0_25), .ZN(n_2_700));
   NOR2_X1 i_2_0_882 (.A1(n_2_0_56), .A2(n_2_0_26), .ZN(n_2_701));
   NOR2_X1 i_2_0_883 (.A1(n_2_0_56), .A2(n_2_0_27), .ZN(n_2_702));
   NOR2_X1 i_2_0_884 (.A1(n_2_0_56), .A2(n_2_0_28), .ZN(n_2_712));
   NOR2_X1 i_2_0_885 (.A1(n_2_0_56), .A2(n_2_0_29), .ZN(n_2_713__0));
   NOR2_X1 i_2_0_886 (.A1(n_2_0_56), .A2(n_2_0_30), .ZN(n_2_714__0));
   NOR2_X1 i_2_0_887 (.A1(n_2_0_56), .A2(n_2_0_31), .ZN(n_2_779));
   NOR2_X1 i_2_0_888 (.A1(n_2_0_56), .A2(n_2_0_32), .ZN(n_2_846));
   INV_X1 i_2_0_889 (.A(n_793), .ZN(n_2_0_57));
   NOR2_X1 i_2_0_890 (.A1(n_2_0_57), .A2(n_2_0_1), .ZN(n_165));
   NOR2_X1 i_2_0_891 (.A1(n_2_0_57), .A2(n_2_0_2), .ZN(n_166));
   NOR2_X1 i_2_0_892 (.A1(n_2_0_57), .A2(n_2_0_3), .ZN(n_167));
   NOR2_X1 i_2_0_893 (.A1(n_2_0_57), .A2(n_2_0_4), .ZN(n_168));
   NOR2_X1 i_2_0_894 (.A1(n_2_0_57), .A2(n_2_0_5), .ZN(n_169));
   NOR2_X1 i_2_0_895 (.A1(n_2_0_57), .A2(n_2_0_6), .ZN(n_170));
   NOR2_X1 i_2_0_896 (.A1(n_2_0_57), .A2(n_2_0_7), .ZN(n_171));
   NOR2_X1 i_2_0_897 (.A1(n_2_0_57), .A2(n_2_0_8), .ZN(n_172));
   NOR2_X1 i_2_0_898 (.A1(n_2_0_57), .A2(n_2_0_9), .ZN(n_173));
   NOR2_X1 i_2_0_899 (.A1(n_2_0_57), .A2(n_2_0_10), .ZN(n_174));
   NOR2_X1 i_2_0_900 (.A1(n_2_0_57), .A2(n_2_0_11), .ZN(n_175));
   NOR2_X1 i_2_0_901 (.A1(n_2_0_57), .A2(n_2_0_12), .ZN(n_176));
   NOR2_X1 i_2_0_902 (.A1(n_2_0_57), .A2(n_2_0_13), .ZN(n_177));
   NOR2_X1 i_2_0_903 (.A1(n_2_0_57), .A2(n_2_0_14), .ZN(n_178));
   NOR2_X1 i_2_0_904 (.A1(n_2_0_57), .A2(n_2_0_15), .ZN(n_179));
   NOR2_X1 i_2_0_905 (.A1(n_2_0_57), .A2(n_2_0_16), .ZN(n_180));
   NOR2_X1 i_2_0_906 (.A1(n_2_0_57), .A2(n_2_0_17), .ZN(n_181));
   NOR2_X1 i_2_0_907 (.A1(n_2_0_57), .A2(n_2_0_18), .ZN(n_182));
   NOR2_X1 i_2_0_908 (.A1(n_2_0_57), .A2(n_2_0_19), .ZN(n_183));
   NOR2_X1 i_2_0_909 (.A1(n_2_0_57), .A2(n_2_0_20), .ZN(n_184));
   NOR2_X1 i_2_0_910 (.A1(n_2_0_57), .A2(n_2_0_21), .ZN(n_185));
   NOR2_X1 i_2_0_911 (.A1(n_2_0_57), .A2(n_2_0_22), .ZN(n_186));
   NOR2_X1 i_2_0_912 (.A1(n_2_0_57), .A2(n_2_0_23), .ZN(n_187));
   NOR2_X1 i_2_0_913 (.A1(n_2_0_57), .A2(n_2_0_24), .ZN(n_188));
   NOR2_X1 i_2_0_914 (.A1(n_2_0_57), .A2(n_2_0_25), .ZN(n_189));
   NOR2_X1 i_2_0_915 (.A1(n_2_0_57), .A2(n_2_0_26), .ZN(n_190));
   NOR2_X1 i_2_0_916 (.A1(n_2_0_57), .A2(n_2_0_27), .ZN(n_191));
   NOR2_X1 i_2_0_917 (.A1(n_2_0_57), .A2(n_2_0_28), .ZN(n_192));
   NOR2_X1 i_2_0_918 (.A1(n_2_0_57), .A2(n_2_0_29), .ZN(n_193));
   NOR2_X1 i_2_0_919 (.A1(n_2_0_57), .A2(n_2_0_30), .ZN(n_194));
   NOR2_X1 i_2_0_920 (.A1(n_2_0_57), .A2(n_2_0_31), .ZN(n_195));
   NOR2_X1 i_2_0_921 (.A1(n_2_0_57), .A2(n_2_0_32), .ZN(n_196));
   INV_X1 i_2_0_922 (.A(n_792), .ZN(n_2_0_58));
   NOR2_X1 i_2_0_923 (.A1(n_2_0_58), .A2(n_2_0_1), .ZN(n_197));
   NOR2_X1 i_2_0_924 (.A1(n_2_0_58), .A2(n_2_0_2), .ZN(n_198));
   NOR2_X1 i_2_0_925 (.A1(n_2_0_58), .A2(n_2_0_3), .ZN(n_199));
   NOR2_X1 i_2_0_926 (.A1(n_2_0_58), .A2(n_2_0_4), .ZN(n_200));
   NOR2_X1 i_2_0_927 (.A1(n_2_0_58), .A2(n_2_0_5), .ZN(n_201));
   NOR2_X1 i_2_0_928 (.A1(n_2_0_58), .A2(n_2_0_6), .ZN(n_202));
   NOR2_X1 i_2_0_929 (.A1(n_2_0_58), .A2(n_2_0_7), .ZN(n_203));
   NOR2_X1 i_2_0_930 (.A1(n_2_0_58), .A2(n_2_0_8), .ZN(n_204));
   NOR2_X1 i_2_0_931 (.A1(n_2_0_58), .A2(n_2_0_9), .ZN(n_205));
   NOR2_X1 i_2_0_932 (.A1(n_2_0_58), .A2(n_2_0_10), .ZN(n_206));
   NOR2_X1 i_2_0_933 (.A1(n_2_0_58), .A2(n_2_0_11), .ZN(n_207));
   NOR2_X1 i_2_0_934 (.A1(n_2_0_58), .A2(n_2_0_12), .ZN(n_208));
   NOR2_X1 i_2_0_935 (.A1(n_2_0_58), .A2(n_2_0_13), .ZN(n_209));
   NOR2_X1 i_2_0_936 (.A1(n_2_0_58), .A2(n_2_0_14), .ZN(n_210));
   NOR2_X1 i_2_0_937 (.A1(n_2_0_58), .A2(n_2_0_15), .ZN(n_211));
   NOR2_X1 i_2_0_938 (.A1(n_2_0_58), .A2(n_2_0_16), .ZN(n_212));
   NOR2_X1 i_2_0_939 (.A1(n_2_0_58), .A2(n_2_0_17), .ZN(n_213));
   NOR2_X1 i_2_0_940 (.A1(n_2_0_58), .A2(n_2_0_18), .ZN(n_214));
   NOR2_X1 i_2_0_941 (.A1(n_2_0_58), .A2(n_2_0_19), .ZN(n_215));
   NOR2_X1 i_2_0_942 (.A1(n_2_0_58), .A2(n_2_0_20), .ZN(n_216));
   NOR2_X1 i_2_0_943 (.A1(n_2_0_58), .A2(n_2_0_21), .ZN(n_217));
   NOR2_X1 i_2_0_944 (.A1(n_2_0_58), .A2(n_2_0_22), .ZN(n_218));
   NOR2_X1 i_2_0_945 (.A1(n_2_0_58), .A2(n_2_0_23), .ZN(n_219));
   NOR2_X1 i_2_0_946 (.A1(n_2_0_58), .A2(n_2_0_24), .ZN(n_220));
   NOR2_X1 i_2_0_947 (.A1(n_2_0_58), .A2(n_2_0_25), .ZN(n_221));
   NOR2_X1 i_2_0_948 (.A1(n_2_0_58), .A2(n_2_0_26), .ZN(n_222));
   NOR2_X1 i_2_0_949 (.A1(n_2_0_58), .A2(n_2_0_27), .ZN(n_223));
   NOR2_X1 i_2_0_950 (.A1(n_2_0_58), .A2(n_2_0_28), .ZN(n_224));
   NOR2_X1 i_2_0_951 (.A1(n_2_0_58), .A2(n_2_0_29), .ZN(n_225));
   NOR2_X1 i_2_0_952 (.A1(n_2_0_58), .A2(n_2_0_30), .ZN(n_226));
   NOR2_X1 i_2_0_953 (.A1(n_2_0_58), .A2(n_2_0_31), .ZN(n_227));
   NOR2_X1 i_2_0_954 (.A1(n_2_0_58), .A2(n_2_0_32), .ZN(n_228));
   INV_X1 i_2_0_955 (.A(n_791), .ZN(n_2_0_59));
   NOR2_X1 i_2_0_956 (.A1(n_2_0_59), .A2(n_2_0_1), .ZN(n_229));
   NOR2_X1 i_2_0_957 (.A1(n_2_0_59), .A2(n_2_0_2), .ZN(n_230));
   NOR2_X1 i_2_0_958 (.A1(n_2_0_59), .A2(n_2_0_3), .ZN(n_231));
   NOR2_X1 i_2_0_959 (.A1(n_2_0_59), .A2(n_2_0_4), .ZN(n_232));
   NOR2_X1 i_2_0_960 (.A1(n_2_0_59), .A2(n_2_0_5), .ZN(n_233));
   NOR2_X1 i_2_0_961 (.A1(n_2_0_59), .A2(n_2_0_6), .ZN(n_234));
   NOR2_X1 i_2_0_962 (.A1(n_2_0_59), .A2(n_2_0_7), .ZN(n_235));
   NOR2_X1 i_2_0_963 (.A1(n_2_0_59), .A2(n_2_0_8), .ZN(n_236));
   NOR2_X1 i_2_0_964 (.A1(n_2_0_59), .A2(n_2_0_9), .ZN(n_237));
   NOR2_X1 i_2_0_965 (.A1(n_2_0_59), .A2(n_2_0_10), .ZN(n_238));
   NOR2_X1 i_2_0_966 (.A1(n_2_0_59), .A2(n_2_0_11), .ZN(n_239));
   NOR2_X1 i_2_0_967 (.A1(n_2_0_59), .A2(n_2_0_12), .ZN(n_240));
   NOR2_X1 i_2_0_968 (.A1(n_2_0_59), .A2(n_2_0_13), .ZN(n_241));
   NOR2_X1 i_2_0_969 (.A1(n_2_0_59), .A2(n_2_0_14), .ZN(n_242));
   NOR2_X1 i_2_0_970 (.A1(n_2_0_59), .A2(n_2_0_15), .ZN(n_243));
   NOR2_X1 i_2_0_971 (.A1(n_2_0_59), .A2(n_2_0_16), .ZN(n_244));
   NOR2_X1 i_2_0_972 (.A1(n_2_0_59), .A2(n_2_0_17), .ZN(n_245));
   NOR2_X1 i_2_0_973 (.A1(n_2_0_59), .A2(n_2_0_18), .ZN(n_246));
   NOR2_X1 i_2_0_974 (.A1(n_2_0_59), .A2(n_2_0_19), .ZN(n_247));
   NOR2_X1 i_2_0_975 (.A1(n_2_0_59), .A2(n_2_0_20), .ZN(n_248));
   NOR2_X1 i_2_0_976 (.A1(n_2_0_59), .A2(n_2_0_21), .ZN(n_249));
   NOR2_X1 i_2_0_977 (.A1(n_2_0_59), .A2(n_2_0_22), .ZN(n_250));
   NOR2_X1 i_2_0_978 (.A1(n_2_0_59), .A2(n_2_0_23), .ZN(n_251));
   NOR2_X1 i_2_0_979 (.A1(n_2_0_59), .A2(n_2_0_24), .ZN(n_252));
   NOR2_X1 i_2_0_980 (.A1(n_2_0_59), .A2(n_2_0_25), .ZN(n_253));
   NOR2_X1 i_2_0_981 (.A1(n_2_0_59), .A2(n_2_0_26), .ZN(n_254));
   NOR2_X1 i_2_0_982 (.A1(n_2_0_59), .A2(n_2_0_27), .ZN(n_255));
   NOR2_X1 i_2_0_983 (.A1(n_2_0_59), .A2(n_2_0_28), .ZN(n_256));
   NOR2_X1 i_2_0_984 (.A1(n_2_0_59), .A2(n_2_0_29), .ZN(n_257));
   NOR2_X1 i_2_0_985 (.A1(n_2_0_59), .A2(n_2_0_30), .ZN(n_258));
   NOR2_X1 i_2_0_986 (.A1(n_2_0_59), .A2(n_2_0_31), .ZN(n_259));
   NOR2_X1 i_2_0_987 (.A1(n_2_0_59), .A2(n_2_0_32), .ZN(n_260));
   INV_X1 i_2_0_988 (.A(n_790), .ZN(n_2_0_60));
   NOR2_X1 i_2_0_989 (.A1(n_2_0_60), .A2(n_2_0_1), .ZN(n_261));
   NOR2_X1 i_2_0_990 (.A1(n_2_0_60), .A2(n_2_0_2), .ZN(n_262));
   NOR2_X1 i_2_0_991 (.A1(n_2_0_60), .A2(n_2_0_3), .ZN(n_263));
   NOR2_X1 i_2_0_992 (.A1(n_2_0_60), .A2(n_2_0_4), .ZN(n_264));
   NOR2_X1 i_2_0_993 (.A1(n_2_0_60), .A2(n_2_0_5), .ZN(n_265));
   NOR2_X1 i_2_0_994 (.A1(n_2_0_60), .A2(n_2_0_6), .ZN(n_266));
   NOR2_X1 i_2_0_995 (.A1(n_2_0_60), .A2(n_2_0_7), .ZN(n_267));
   NOR2_X1 i_2_0_996 (.A1(n_2_0_60), .A2(n_2_0_8), .ZN(n_268));
   NOR2_X1 i_2_0_997 (.A1(n_2_0_60), .A2(n_2_0_9), .ZN(n_269));
   NOR2_X1 i_2_0_998 (.A1(n_2_0_60), .A2(n_2_0_10), .ZN(n_270));
   NOR2_X1 i_2_0_999 (.A1(n_2_0_60), .A2(n_2_0_11), .ZN(n_271));
   NOR2_X1 i_2_0_1000 (.A1(n_2_0_60), .A2(n_2_0_12), .ZN(n_272));
   NOR2_X1 i_2_0_1001 (.A1(n_2_0_60), .A2(n_2_0_13), .ZN(n_273));
   NOR2_X1 i_2_0_1002 (.A1(n_2_0_60), .A2(n_2_0_14), .ZN(n_274));
   NOR2_X1 i_2_0_1003 (.A1(n_2_0_60), .A2(n_2_0_15), .ZN(n_275));
   NOR2_X1 i_2_0_1004 (.A1(n_2_0_60), .A2(n_2_0_16), .ZN(n_276));
   NOR2_X1 i_2_0_1005 (.A1(n_2_0_60), .A2(n_2_0_17), .ZN(n_277));
   NOR2_X1 i_2_0_1006 (.A1(n_2_0_60), .A2(n_2_0_18), .ZN(n_278));
   NOR2_X1 i_2_0_1007 (.A1(n_2_0_60), .A2(n_2_0_19), .ZN(n_279));
   NOR2_X1 i_2_0_1008 (.A1(n_2_0_60), .A2(n_2_0_20), .ZN(n_280));
   NOR2_X1 i_2_0_1009 (.A1(n_2_0_60), .A2(n_2_0_21), .ZN(n_281));
   NOR2_X1 i_2_0_1010 (.A1(n_2_0_60), .A2(n_2_0_22), .ZN(n_282));
   NOR2_X1 i_2_0_1011 (.A1(n_2_0_60), .A2(n_2_0_23), .ZN(n_283));
   NOR2_X1 i_2_0_1012 (.A1(n_2_0_60), .A2(n_2_0_24), .ZN(n_284));
   NOR2_X1 i_2_0_1013 (.A1(n_2_0_60), .A2(n_2_0_25), .ZN(n_285));
   NOR2_X1 i_2_0_1014 (.A1(n_2_0_60), .A2(n_2_0_26), .ZN(n_286));
   NOR2_X1 i_2_0_1015 (.A1(n_2_0_60), .A2(n_2_0_27), .ZN(n_287));
   NOR2_X1 i_2_0_1016 (.A1(n_2_0_60), .A2(n_2_0_28), .ZN(n_288));
   NOR2_X1 i_2_0_1017 (.A1(n_2_0_60), .A2(n_2_0_29), .ZN(n_289));
   NOR2_X1 i_2_0_1018 (.A1(n_2_0_60), .A2(n_2_0_30), .ZN(n_290));
   NOR2_X1 i_2_0_1019 (.A1(n_2_0_60), .A2(n_2_0_31), .ZN(n_291));
   NOR2_X1 i_2_0_1020 (.A1(n_2_0_60), .A2(n_2_0_32), .ZN(n_292));
   INV_X1 i_2_0_1021 (.A(n_789), .ZN(n_2_0_61));
   NOR2_X1 i_2_0_1022 (.A1(n_2_0_61), .A2(n_2_0_1), .ZN(n_293));
   NOR2_X1 i_2_0_1023 (.A1(n_2_0_61), .A2(n_2_0_2), .ZN(n_294));
   NOR2_X1 i_2_0_1024 (.A1(n_2_0_61), .A2(n_2_0_3), .ZN(n_295));
   NOR2_X1 i_2_0_1025 (.A1(n_2_0_61), .A2(n_2_0_4), .ZN(n_296));
   NOR2_X1 i_2_0_1026 (.A1(n_2_0_61), .A2(n_2_0_5), .ZN(n_297));
   NOR2_X1 i_2_0_1027 (.A1(n_2_0_61), .A2(n_2_0_6), .ZN(n_298));
   NOR2_X1 i_2_0_1028 (.A1(n_2_0_61), .A2(n_2_0_7), .ZN(n_299));
   NOR2_X1 i_2_0_1029 (.A1(n_2_0_61), .A2(n_2_0_8), .ZN(n_300));
   NOR2_X1 i_2_0_1030 (.A1(n_2_0_61), .A2(n_2_0_9), .ZN(n_301));
   NOR2_X1 i_2_0_1031 (.A1(n_2_0_61), .A2(n_2_0_10), .ZN(n_302));
   NOR2_X1 i_2_0_1032 (.A1(n_2_0_61), .A2(n_2_0_11), .ZN(n_303));
   NOR2_X1 i_2_0_1033 (.A1(n_2_0_61), .A2(n_2_0_12), .ZN(n_304));
   NOR2_X1 i_2_0_1034 (.A1(n_2_0_61), .A2(n_2_0_13), .ZN(n_305));
   NOR2_X1 i_2_0_1035 (.A1(n_2_0_61), .A2(n_2_0_14), .ZN(n_306));
   NOR2_X1 i_2_0_1036 (.A1(n_2_0_61), .A2(n_2_0_15), .ZN(n_307));
   NOR2_X1 i_2_0_1037 (.A1(n_2_0_61), .A2(n_2_0_16), .ZN(n_308));
   NOR2_X1 i_2_0_1038 (.A1(n_2_0_61), .A2(n_2_0_17), .ZN(n_309));
   NOR2_X1 i_2_0_1039 (.A1(n_2_0_61), .A2(n_2_0_18), .ZN(n_310));
   NOR2_X1 i_2_0_1040 (.A1(n_2_0_61), .A2(n_2_0_19), .ZN(n_311));
   NOR2_X1 i_2_0_1041 (.A1(n_2_0_61), .A2(n_2_0_20), .ZN(n_312));
   NOR2_X1 i_2_0_1042 (.A1(n_2_0_61), .A2(n_2_0_21), .ZN(n_313));
   NOR2_X1 i_2_0_1043 (.A1(n_2_0_61), .A2(n_2_0_22), .ZN(n_314));
   NOR2_X1 i_2_0_1044 (.A1(n_2_0_61), .A2(n_2_0_23), .ZN(n_315));
   NOR2_X1 i_2_0_1045 (.A1(n_2_0_61), .A2(n_2_0_24), .ZN(n_316));
   NOR2_X1 i_2_0_1046 (.A1(n_2_0_61), .A2(n_2_0_25), .ZN(n_317));
   NOR2_X1 i_2_0_1047 (.A1(n_2_0_61), .A2(n_2_0_26), .ZN(n_318));
   NOR2_X1 i_2_0_1048 (.A1(n_2_0_61), .A2(n_2_0_27), .ZN(n_319));
   NOR2_X1 i_2_0_1049 (.A1(n_2_0_61), .A2(n_2_0_28), .ZN(n_320));
   NOR2_X1 i_2_0_1050 (.A1(n_2_0_61), .A2(n_2_0_29), .ZN(n_321));
   NOR2_X1 i_2_0_1051 (.A1(n_2_0_61), .A2(n_2_0_30), .ZN(n_322));
   NOR2_X1 i_2_0_1052 (.A1(n_2_0_61), .A2(n_2_0_31), .ZN(n_323));
   NOR2_X1 i_2_0_1053 (.A1(n_2_0_61), .A2(n_2_0_32), .ZN(n_324));
   INV_X1 i_2_0_1054 (.A(y), .ZN(n_2_0_62));
   NOR2_X1 i_2_0_1055 (.A1(n_2_0_1), .A2(n_2_0_62), .ZN(n_325));
   NOR2_X1 i_2_0_1056 (.A1(n_2_0_2), .A2(n_2_0_62), .ZN(n_326));
   NOR2_X1 i_2_0_1057 (.A1(n_2_0_3), .A2(n_2_0_62), .ZN(n_327));
   NOR2_X1 i_2_0_1058 (.A1(n_2_0_4), .A2(n_2_0_62), .ZN(n_328));
   NOR2_X1 i_2_0_1059 (.A1(n_2_0_5), .A2(n_2_0_62), .ZN(n_329));
   NOR2_X1 i_2_0_1060 (.A1(n_2_0_6), .A2(n_2_0_62), .ZN(n_330));
   NOR2_X1 i_2_0_1061 (.A1(n_2_0_7), .A2(n_2_0_62), .ZN(n_331));
   NOR2_X1 i_2_0_1062 (.A1(n_2_0_8), .A2(n_2_0_62), .ZN(n_332));
   NOR2_X1 i_2_0_1063 (.A1(n_2_0_9), .A2(n_2_0_62), .ZN(n_333));
   NOR2_X1 i_2_0_1064 (.A1(n_2_0_10), .A2(n_2_0_62), .ZN(n_334));
   NOR2_X1 i_2_0_1065 (.A1(n_2_0_11), .A2(n_2_0_62), .ZN(n_335));
   NOR2_X1 i_2_0_1066 (.A1(n_2_0_12), .A2(n_2_0_62), .ZN(n_336));
   NOR2_X1 i_2_0_1067 (.A1(n_2_0_13), .A2(n_2_0_62), .ZN(n_337));
   NOR2_X1 i_2_0_1068 (.A1(n_2_0_14), .A2(n_2_0_62), .ZN(n_338));
   NOR2_X1 i_2_0_1069 (.A1(n_2_0_15), .A2(n_2_0_62), .ZN(n_339));
   NOR2_X1 i_2_0_1070 (.A1(n_2_0_16), .A2(n_2_0_62), .ZN(n_340));
   NOR2_X1 i_2_0_1071 (.A1(n_2_0_17), .A2(n_2_0_62), .ZN(n_341));
   NOR2_X1 i_2_0_1072 (.A1(n_2_0_18), .A2(n_2_0_62), .ZN(n_342));
   NOR2_X1 i_2_0_1073 (.A1(n_2_0_19), .A2(n_2_0_62), .ZN(n_343));
   NOR2_X1 i_2_0_1074 (.A1(n_2_0_20), .A2(n_2_0_62), .ZN(n_344));
   NOR2_X1 i_2_0_1075 (.A1(n_2_0_21), .A2(n_2_0_62), .ZN(n_345));
   NOR2_X1 i_2_0_1076 (.A1(n_2_0_22), .A2(n_2_0_62), .ZN(n_346));
   NOR2_X1 i_2_0_1077 (.A1(n_2_0_23), .A2(n_2_0_62), .ZN(n_347));
   NOR2_X1 i_2_0_1078 (.A1(n_2_0_24), .A2(n_2_0_62), .ZN(n_348));
   NOR2_X1 i_2_0_1079 (.A1(n_2_0_25), .A2(n_2_0_62), .ZN(n_349));
   NOR2_X1 i_2_0_1080 (.A1(n_2_0_26), .A2(n_2_0_62), .ZN(n_350));
   NOR2_X1 i_2_0_1081 (.A1(n_2_0_27), .A2(n_2_0_62), .ZN(n_351));
   NOR2_X1 i_2_0_1082 (.A1(n_2_0_28), .A2(n_2_0_62), .ZN(n_352));
   NOR2_X1 i_2_0_1083 (.A1(n_2_0_29), .A2(n_2_0_62), .ZN(n_353));
   NOR2_X1 i_2_0_1084 (.A1(n_2_0_30), .A2(n_2_0_62), .ZN(n_354));
   NOR2_X1 i_2_0_1085 (.A1(n_2_0_31), .A2(n_2_0_62), .ZN(n_355));
   NOR2_X1 i_2_0_1086 (.A1(n_2_0_32), .A2(n_2_0_62), .ZN(n_356));
   CSA__1_2043 cs6 (.x({n_2_643, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, 
      uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, n_2_642, n_2_641, n_2_640, 
      n_2_639, n_2_638, n_2_637, n_2_636, n_2_635, n_2_634, n_2_633, n_2_632, 
      n_2_631, n_2_630, n_2_629, n_2_628, n_2_627, n_2_626, n_2_625, n_2_624, 
      n_2_623, n_2_622, n_2_621, n_2_620, n_2_619, n_2_618, n_2_617, n_2_616, 
      n_2_615, n_2_614, n_2_613, uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, 
      uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, 
      uc_64, uc_65}), .y({n_2_675, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, 
      uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, n_2_674, n_2_673, n_2_672, 
      n_2_671, n_2_670, n_2_669, n_2_668, n_2_667, n_2_666, n_2_665, n_2_664, 
      n_2_663, n_2_662, n_2_661, n_2_660, n_2_659, n_2_658, n_2_657, n_2_656, 
      n_2_655, n_2_654, n_2_653, n_2_652, n_2_651, n_2_650, n_2_649, n_2_648, 
      n_2_647, n_2_646, n_2_645, n_2_644, uc_79, uc_80, uc_81, uc_82, uc_83, 
      uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, 
      uc_94, uc_95, uc_96, uc_97}), .z({n_2_846, uc_98, uc_99, uc_100, uc_101, 
      uc_102, uc_103, uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, n_2_779, 
      n_2_714__0, n_2_713__0, n_2_712, n_2_702, n_2_701, n_2_700, n_2_699, 
      n_2_698, n_2_697, n_2_696, n_2_695, n_2_694, n_2_693, n_2_692, n_2_691, 
      n_2_690, n_2_689, n_2_688, n_2_687, n_2_686, n_2_685, n_2_684, n_2_683, 
      n_2_682, n_2_681, n_2_680, n_2_679, n_2_678, n_2_677, n_2_676, uc_110, 
      uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, uc_118, uc_119, 
      uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, uc_126, uc_127, uc_128, 
      uc_129}), .s({n_401, n_400, n_399, n_398, n_397, n_396, n_395, n_394, 
      n_393, n_392, n_391, n_390, n_389, n_388, n_387, n_386, n_385, n_384, 
      n_383, n_382, n_381, n_380, n_379, n_378, n_377, n_376, n_375, n_374, 
      n_373, n_372, n_371, n_370, n_369, n_368, n_367, n_366, n_365, n_364, 
      n_363, n_362, n_361, n_360, n_359, n_358, n_357, uc_130, uc_131, uc_132, 
      uc_133, uc_134, uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, 
      uc_142, uc_143, uc_144, uc_145, uc_146, uc_147, uc_148}), .carry_final());
   CSA__1_3068 cs0 (.x({n_2_71, uc_149, uc_150, uc_151, uc_152, uc_153, uc_154, 
      uc_155, uc_156, uc_157, uc_158, uc_159, uc_160, uc_161, uc_162, uc_163, 
      uc_164, uc_165, uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, uc_172, 
      uc_173, uc_174, uc_175, uc_176, uc_177, uc_178, uc_179, uc_180, n_2_70, 
      n_2_69, n_2_68, n_2_67, n_2_66, n_2_65, n_2_64, n_2_63, n_2_62, n_2_61, 
      n_2_60, n_2_59, n_2_58, n_2_57, n_2_56, n_2_55, n_2_54, n_2_53, n_2_52, 
      n_2_51, n_2_50, n_2_49, n_2_48, n_2_47, n_2_46, n_2_45, n_2_44, n_2_43, 
      n_2_42, n_2_41, uc_181}), .y({n_2_103, uc_182, uc_183, uc_184, uc_185, 
      uc_186, uc_187, uc_188, uc_189, uc_190, uc_191, uc_192, uc_193, uc_194, 
      uc_195, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, 
      uc_204, uc_205, uc_206, uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, 
      n_2_102, n_2_101, n_2_100, n_2_99, n_2_98, n_2_97, n_2_96, n_2_95, n_2_94, 
      n_2_93, n_2_92, n_2_91, n_2_90, n_2_89, n_2_88, n_2_87, n_2_86, n_2_85, 
      n_2_84, n_2_83, n_2_82, n_2_81, n_2_80, n_2_79, n_2_78, n_2_77, n_2_76, 
      n_2_75, n_2_74, n_2_73, n_2_72, uc_213}), .z({n_2_135, uc_214, uc_215, 
      uc_216, uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, uc_223, uc_224, 
      uc_225, uc_226, uc_227, uc_228, uc_229, uc_230, uc_231, uc_232, uc_233, 
      uc_234, uc_235, uc_236, uc_237, uc_238, uc_239, uc_240, uc_241, uc_242, 
      uc_243, n_2_134, n_2_133, n_2_132, n_2_131, n_2_130, n_2_129, n_2_128, 
      n_2_127, n_2_126, n_2_125, n_2_124, n_2_123, n_2_122, n_2_121, n_2_120, 
      n_2_119, n_2_118, n_2_117, n_2_116, n_2_115, n_2_114, n_2_113, n_2_112, 
      n_2_111, n_2_110, n_2_109, n_2_108, n_2_107, n_2_106, n_2_105, n_2_104, 
      uc_244, uc_245}), .s({n_464, n_463, n_462, n_461, n_460, n_459, n_458, 
      n_457, n_456, n_455, n_454, n_453, n_452, n_451, n_450, n_449, n_448, 
      n_447, n_446, n_445, n_444, n_443, n_442, n_441, n_440, n_439, n_438, 
      n_437, n_436, n_435, n_434, n_433, n_432, n_431, n_430, n_429, n_428, 
      n_427, n_426, n_425, n_424, n_423, n_422, n_421, n_420, n_419, n_418, 
      n_417, n_416, n_415, n_414, n_413, n_412, n_411, n_410, n_409, n_408, 
      n_407, n_406, n_405, n_404, n_403, n_402, uc_246}), .carry_final());
   CSA__1_4093 cs1 (.x({n_2_166, uc_247, uc_248, uc_249, uc_250, uc_251, uc_252, 
      uc_253, uc_254, uc_255, uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, 
      uc_262, uc_263, uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, 
      uc_271, uc_272, uc_273, uc_274, uc_275, n_2_165, n_2_164, n_2_163, n_2_162, 
      n_2_161, n_2_160, n_2_159, n_2_158, n_2_157, n_2_156, n_2_155, n_2_154, 
      n_2_153, n_2_152, n_2_151, n_2_150, n_2_149, n_2_148, n_2_147, n_2_146, 
      n_2_145, n_2_144, n_2_143, n_2_142, n_2_141, n_2_140, n_2_139, n_2_138, 
      n_2_137, n_2_136, uc_276, uc_277, uc_278, uc_279}), .y({n_2_198, uc_280, 
      uc_281, uc_282, uc_283, uc_284, uc_285, uc_286, uc_287, uc_288, uc_289, 
      uc_290, uc_291, uc_292, uc_293, uc_294, uc_295, uc_296, uc_297, uc_298, 
      uc_299, uc_300, uc_301, uc_302, uc_303, uc_304, uc_305, uc_306, uc_307, 
      n_2_197, n_2_196, n_2_195, n_2_194, n_2_193, n_2_192, n_2_191, n_2_190, 
      n_2_189, n_2_188, n_2_187, n_2_186, n_2_185, n_2_184, n_2_183, n_2_182, 
      n_2_181, n_2_180, n_2_179, n_2_178, n_2_177, n_2_176, n_2_175, n_2_174, 
      n_2_173, n_2_172, n_2_171, n_2_170, n_2_169, n_2_168, n_2_167, uc_308, 
      uc_309, uc_310, uc_311}), .z({n_2_230, uc_312, uc_313, uc_314, uc_315, 
      uc_316, uc_317, uc_318, uc_319, uc_320, uc_321, uc_322, uc_323, uc_324, 
      uc_325, uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, 
      uc_334, uc_335, uc_336, uc_337, uc_338, n_2_229, n_2_228, n_2_227, n_2_226, 
      n_2_225, n_2_224, n_2_223, n_2_222, n_2_221, n_2_220, n_2_219, n_2_218, 
      n_2_217, n_2_216, n_2_215, n_2_214, n_2_213, n_2_212, n_2_211, n_2_210, 
      n_2_209, n_2_208, n_2_207, n_2_206, n_2_205, n_2_204, n_2_203, n_2_202, 
      n_2_201, n_2_200, n_2_199, uc_339, uc_340, uc_341, uc_342, uc_343}), 
      .s({n_524, n_523, n_522, n_521, n_520, n_519, n_518, n_517, n_516, n_515, 
      n_514, n_513, n_512, n_511, n_510, n_509, n_508, n_507, n_506, n_505, 
      n_504, n_503, n_502, n_501, n_500, n_499, n_498, n_497, n_496, n_495, 
      n_494, n_493, n_492, n_491, n_490, n_489, n_488, n_487, n_486, n_485, 
      n_484, n_483, n_482, n_481, n_480, n_479, n_478, n_477, n_476, n_475, 
      n_474, n_473, n_472, n_471, n_470, n_469, n_468, n_467, n_466, n_465, 
      uc_344, uc_345, uc_346, uc_347}), .carry_final());
   CSA__1_5118 cs2 (.x({n_2_261, uc_348, uc_349, uc_350, uc_351, uc_352, uc_353, 
      uc_354, uc_355, uc_356, uc_357, uc_358, uc_359, uc_360, uc_361, uc_362, 
      uc_363, uc_364, uc_365, uc_366, uc_367, uc_368, uc_369, uc_370, uc_371, 
      uc_372, uc_373, n_2_260, n_2_259, n_2_258, n_2_257, n_2_256, n_2_255, 
      n_2_254, n_2_253, n_2_252, n_2_251, n_2_250, n_2_249, n_2_248, n_2_247, 
      n_2_246, n_2_245, n_2_244, n_2_243, n_2_242, n_2_241, n_2_240, n_2_239, 
      n_2_238, n_2_237, n_2_236, n_2_235, n_2_234, n_2_233, n_2_232, n_2_231, 
      uc_374, uc_375, uc_376, uc_377, uc_378, uc_379, uc_380}), .y({n_2_293, 
      uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, uc_389, 
      uc_390, uc_391, uc_392, uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, 
      uc_399, uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, n_2_292, n_2_291, 
      n_2_290, n_2_289, n_2_288, n_2_287, n_2_286, n_2_285, n_2_284, n_2_283, 
      n_2_282, n_2_281, n_2_280, n_2_279, n_2_278, n_2_277, n_2_276, n_2_275, 
      n_2_274, n_2_273, n_2_272, n_2_271, n_2_270, n_2_269, n_2_268, n_2_267, 
      n_2_266, n_2_265, n_2_264, n_2_263, n_2_262, uc_406, uc_407, uc_408, 
      uc_409, uc_410, uc_411, uc_412}), .z({n_2_325, uc_413, uc_414, uc_415, 
      uc_416, uc_417, uc_418, uc_419, uc_420, uc_421, uc_422, uc_423, uc_424, 
      uc_425, uc_426, uc_427, uc_428, uc_429, uc_430, uc_431, uc_432, uc_433, 
      uc_434, uc_435, uc_436, n_2_324, n_2_323, n_2_322, n_2_321, n_2_320, 
      n_2_319, n_2_318, n_2_317, n_2_316, n_2_315, n_2_314, n_2_313, n_2_312, 
      n_2_311, n_2_310, n_2_309, n_2_308, n_2_307, n_2_306, n_2_305, n_2_304, 
      n_2_303, n_2_302, n_2_301, n_2_300, n_2_299, n_2_298, n_2_297, n_2_296, 
      n_2_295, n_2_294, uc_437, uc_438, uc_439, uc_440, uc_441, uc_442, uc_443, 
      uc_444}), .s({n_581, n_580, n_579, n_578, n_577, n_576, n_575, n_574, 
      n_573, n_572, n_571, n_570, n_569, n_568, n_567, n_566, n_565, n_564, 
      n_563, n_562, n_561, n_560, n_559, n_558, n_557, n_556, n_555, n_554, 
      n_553, n_552, n_551, n_550, n_549, n_548, n_547, n_546, n_545, n_544, 
      n_543, n_542, n_541, n_540, n_539, n_538, n_537, n_536, n_535, n_534, 
      n_533, n_532, n_531, n_530, n_529, n_528, n_527, n_526, n_525, uc_445, 
      uc_446, uc_447, uc_448, uc_449, uc_450, uc_451}), .carry_final());
   CSA__1_6143 cs11 (.x({n_2_766, n_2_765, n_2_764, n_2_763, n_2_762, n_2_761, 
      n_2_760, n_2_759, n_2_758, n_2_757, n_2_756, n_2_755, n_2_754, n_2_753, 
      n_2_752, n_2_751, n_2_750, n_2_749, n_2_748, n_2_747, n_2_746, n_2_745, 
      n_2_744, n_2_743, n_2_742, n_2_741, n_2_740, n_2_739, n_2_738, n_2_737, 
      n_2_736, n_2_735, n_2_734, n_2_733, n_2_732, n_2_731, n_2_730, n_2_729, 
      n_2_728, n_2_727, n_2_726, n_2_725, n_2_724, n_2_723, n_2_722, n_2_721, 
      n_2_720, n_2_719, n_2_718, n_2_717, n_2_716, n_2_715, uc_452, uc_453, 
      uc_454, uc_455, uc_456, uc_457, uc_458, uc_459, uc_460, uc_461, uc_462, 
      uc_463}), .y({n_2_830, n_2_829, n_2_828, n_2_827, n_2_826, n_2_825, 
      n_2_824, n_2_823, n_2_822, n_2_821, n_2_820, n_2_819, n_2_818, n_2_817, 
      n_2_816, n_2_815, n_2_814, n_2_813, n_2_812, n_2_811, n_2_810, n_2_809, 
      n_2_808, n_2_807, n_2_806, n_2_805, n_2_804, n_2_803, n_2_802, n_2_801, 
      n_2_800, n_2_799, n_2_798, n_2_797, n_2_796, n_2_795, n_2_794, n_2_793, 
      n_2_792, n_2_791, n_2_790, n_2_789, n_2_788, n_2_787, n_2_786, n_2_785, 
      n_2_784, n_2_783, n_2_782, n_2_781, n_2_780, n_2_421, uc_464, uc_465, 
      uc_466, uc_467, uc_468, uc_469, uc_470, uc_471, uc_472, uc_473, uc_474, 
      uc_475}), .z({n_2_845, n_2_844, n_2_843, n_2_842, n_2_841, n_2_840, 
      n_2_839, n_2_838, n_2_837, n_2_836, n_2_835, n_2_834, n_2_833, n_2_832, 
      n_2_831, n_2_778, n_2_777, n_2_776, n_2_775, n_2_774, n_2_773, n_2_772, 
      n_2_771, n_2_770, n_2_769, n_2_768, n_2_767, n_2_711, n_2_710, n_2_709, 
      n_2_708, n_2_707, n_2_706, n_2_705, n_2_704, n_2_703, n_2_9, n_2_8, n_2_7, 
      n_2_6, n_2_5, n_2_4, n_2_3, n_2_2, n_2_1, n_2_0, n_2_848, n_2_847, n_2_517, 
      uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, uc_482, uc_483, uc_484, 
      uc_485, uc_486, uc_487, uc_488, uc_489, uc_490}), .s({n_633, n_632, n_631, 
      n_630, n_629, n_628, n_627, n_626, n_625, n_624, n_623, n_622, n_621, 
      n_620, n_619, n_618, n_617, n_616, n_615, n_614, n_613, n_612, n_611, 
      n_610, n_609, n_608, n_607, n_606, n_605, n_604, n_603, n_602, n_601, 
      n_600, n_599, n_598, n_597, n_596, n_595, n_594, n_593, n_592, n_591, 
      n_590, n_589, n_588, n_587, n_586, n_585, n_584, n_583, n_582, uc_491, 
      uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, uc_499, uc_500, 
      uc_501, uc_502}), .carry_final());
   CSA__1_7168 cs3 (.x({n_2_356, uc_503, uc_504, uc_505, uc_506, uc_507, uc_508, 
      uc_509, uc_510, uc_511, uc_512, uc_513, uc_514, uc_515, uc_516, uc_517, 
      uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, uc_525, n_2_355, 
      n_2_354, n_2_353, n_2_352, n_2_351, n_2_350, n_2_349, n_2_348, n_2_347, 
      n_2_346, n_2_345, n_2_344, n_2_343, n_2_342, n_2_341, n_2_340, n_2_339, 
      n_2_338, n_2_337, n_2_336, n_2_335, n_2_334, n_2_333, n_2_332, n_2_331, 
      n_2_330, n_2_329, n_2_328, n_2_327, n_2_326, uc_526, uc_527, uc_528, 
      uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, uc_535}), .y({n_2_388, 
      uc_536, uc_537, uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, 
      uc_545, uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, 
      uc_554, uc_555, uc_556, uc_557, n_2_387, n_2_386, n_2_385, n_2_384, 
      n_2_383, n_2_382, n_2_381, n_2_380, n_2_379, n_2_378, n_2_377, n_2_376, 
      n_2_375, n_2_374, n_2_373, n_2_372, n_2_371, n_2_370, n_2_369, n_2_368, 
      n_2_367, n_2_366, n_2_365, n_2_364, n_2_363, n_2_362, n_2_361, n_2_360, 
      n_2_359, n_2_358, n_2_357, uc_558, uc_559, uc_560, uc_561, uc_562, uc_563, 
      uc_564, uc_565, uc_566, uc_567}), .z({n_2_420, uc_568, uc_569, uc_570, 
      uc_571, uc_572, uc_573, uc_574, uc_575, uc_576, uc_577, uc_578, uc_579, 
      uc_580, uc_581, uc_582, uc_583, uc_584, uc_585, uc_586, uc_587, uc_588, 
      n_2_419, n_2_418, n_2_417, n_2_416, n_2_415, n_2_414, n_2_413, n_2_412, 
      n_2_411, n_2_410, n_2_409, n_2_408, n_2_407, n_2_406, n_2_405, n_2_404, 
      n_2_403, n_2_402, n_2_401, n_2_400, n_2_399, n_2_398, n_2_397, n_2_396, 
      n_2_395, n_2_394, n_2_393, n_2_392, n_2_391, n_2_390, n_2_389, uc_589, 
      uc_590, uc_591, uc_592, uc_593, uc_594, uc_595, uc_596, uc_597, uc_598, 
      uc_599}), .s({n_2_766, n_2_765, n_2_764, n_2_763, n_2_762, n_2_761, 
      n_2_760, n_2_759, n_2_758, n_2_757, n_2_756, n_2_755, n_2_754, n_2_753, 
      n_2_752, n_2_751, n_2_750, n_2_749, n_2_748, n_2_747, n_2_746, n_2_745, 
      n_2_744, n_2_743, n_2_742, n_2_741, n_2_740, n_2_739, n_2_738, n_2_737, 
      n_2_736, n_2_735, n_2_734, n_2_733, n_2_732, n_2_731, n_2_730, n_2_729, 
      n_2_728, n_2_727, n_2_726, n_2_725, n_2_724, n_2_723, n_2_722, n_2_721, 
      n_2_720, n_2_719, n_2_718, n_2_717, n_2_716, n_2_715, n_2_714__1, 
      n_2_713__1, uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, uc_606, uc_607, 
      uc_608, uc_609}), .carry_final());
   CSA__1_8193 cs4 (.x({n_2_452, uc_610, uc_611, uc_612, uc_613, uc_614, uc_615, 
      uc_616, uc_617, uc_618, uc_619, uc_620, uc_621, uc_622, uc_623, uc_624, 
      uc_625, uc_626, uc_627, uc_628, uc_629, n_2_451, n_2_450, n_2_449, n_2_448, 
      n_2_447, n_2_446, n_2_445, n_2_444, n_2_443, n_2_442, n_2_441, n_2_440, 
      n_2_439, n_2_438, n_2_437, n_2_436, n_2_435, n_2_434, n_2_433, n_2_432, 
      n_2_431, n_2_430, n_2_429, n_2_428, n_2_427, n_2_426, n_2_425, n_2_424, 
      n_2_423, n_2_422, uc_630, uc_631, uc_632, uc_633, uc_634, uc_635, uc_636, 
      uc_637, uc_638, uc_639, uc_640, uc_641, uc_642}), .y({n_2_484, uc_643, 
      uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, uc_651, uc_652, 
      uc_653, uc_654, uc_655, uc_656, uc_657, uc_658, uc_659, uc_660, uc_661, 
      n_2_483, n_2_482, n_2_481, n_2_480, n_2_479, n_2_478, n_2_477, n_2_476, 
      n_2_475, n_2_474, n_2_473, n_2_472, n_2_471, n_2_470, n_2_469, n_2_468, 
      n_2_467, n_2_466, n_2_465, n_2_464, n_2_463, n_2_462, n_2_461, n_2_460, 
      n_2_459, n_2_458, n_2_457, n_2_456, n_2_455, n_2_454, n_2_453, uc_662, 
      uc_663, uc_664, uc_665, uc_666, uc_667, uc_668, uc_669, uc_670, uc_671, 
      uc_672, uc_673, uc_674}), .z({n_2_516, uc_675, uc_676, uc_677, uc_678, 
      uc_679, uc_680, uc_681, uc_682, uc_683, uc_684, uc_685, uc_686, uc_687, 
      uc_688, uc_689, uc_690, uc_691, uc_692, n_2_515, n_2_514, n_2_513, n_2_512, 
      n_2_511, n_2_510, n_2_509, n_2_508, n_2_507, n_2_506, n_2_505, n_2_504, 
      n_2_503, n_2_502, n_2_501, n_2_500, n_2_499, n_2_498, n_2_497, n_2_496, 
      n_2_495, n_2_494, n_2_493, n_2_492, n_2_491, n_2_490, n_2_489, n_2_488, 
      n_2_487, n_2_486, n_2_485, uc_693, uc_694, uc_695, uc_696, uc_697, uc_698, 
      uc_699, uc_700, uc_701, uc_702, uc_703, uc_704, uc_705, uc_706}), .s({
      n_2_830, n_2_829, n_2_828, n_2_827, n_2_826, n_2_825, n_2_824, n_2_823, 
      n_2_822, n_2_821, n_2_820, n_2_819, n_2_818, n_2_817, n_2_816, n_2_815, 
      n_2_814, n_2_813, n_2_812, n_2_811, n_2_810, n_2_809, n_2_808, n_2_807, 
      n_2_806, n_2_805, n_2_804, n_2_803, n_2_802, n_2_801, n_2_800, n_2_799, 
      n_2_798, n_2_797, n_2_796, n_2_795, n_2_794, n_2_793, n_2_792, n_2_791, 
      n_2_790, n_2_789, n_2_788, n_2_787, n_2_786, n_2_785, n_2_784, n_2_783, 
      n_2_782, n_2_781, n_2_780, uc_707, uc_708, uc_709, uc_710, uc_711, uc_712, 
      uc_713, uc_714, uc_715, uc_716, uc_717, uc_718, uc_719}), .carry_final());
   CSA__0_112 cs5 (.x({n_2_548, uc_720, uc_721, uc_722, uc_723, uc_724, uc_725, 
      uc_726, uc_727, uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, uc_734, 
      uc_735, uc_736, n_2_547, n_2_546, n_2_545, n_2_544, n_2_543, n_2_542, 
      n_2_541, n_2_540, n_2_539, n_2_538, n_2_537, n_2_536, n_2_535, n_2_534, 
      n_2_533, n_2_532, n_2_531, n_2_530, n_2_529, n_2_528, n_2_527, n_2_526, 
      n_2_525, n_2_524, n_2_523, n_2_522, n_2_521, n_2_520, n_2_519, n_2_518, 
      uc_737, uc_738, uc_739, uc_740, uc_741, uc_742, uc_743, uc_744, uc_745, 
      uc_746, uc_747, uc_748, uc_749, uc_750, uc_751, uc_752}), .y({n_2_580, 
      uc_753, uc_754, uc_755, uc_756, uc_757, uc_758, uc_759, uc_760, uc_761, 
      uc_762, uc_763, uc_764, uc_765, uc_766, uc_767, uc_768, n_2_579, n_2_578, 
      n_2_577, n_2_576, n_2_575, n_2_574, n_2_573, n_2_572, n_2_571, n_2_570, 
      n_2_569, n_2_568, n_2_567, n_2_566, n_2_565, n_2_564, n_2_563, n_2_562, 
      n_2_561, n_2_560, n_2_559, n_2_558, n_2_557, n_2_556, n_2_555, n_2_554, 
      n_2_553, n_2_552, n_2_551, n_2_550, n_2_549, uc_769, uc_770, uc_771, 
      uc_772, uc_773, uc_774, uc_775, uc_776, uc_777, uc_778, uc_779, uc_780, 
      uc_781, uc_782, uc_783, uc_784}), .z({n_2_612, uc_785, uc_786, uc_787, 
      uc_788, uc_789, uc_790, uc_791, uc_792, uc_793, uc_794, uc_795, uc_796, 
      uc_797, uc_798, uc_799, n_2_611, n_2_610, n_2_609, n_2_608, n_2_607, 
      n_2_606, n_2_605, n_2_604, n_2_603, n_2_602, n_2_601, n_2_600, n_2_599, 
      n_2_598, n_2_597, n_2_596, n_2_595, n_2_594, n_2_593, n_2_592, n_2_591, 
      n_2_590, n_2_589, n_2_588, n_2_587, n_2_586, n_2_585, n_2_584, n_2_583, 
      n_2_582, n_2_581, uc_800, uc_801, uc_802, uc_803, uc_804, uc_805, uc_806, 
      uc_807, uc_808, uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, 
      uc_816}), .s({n_2_845, n_2_844, n_2_843, n_2_842, n_2_841, n_2_840, 
      n_2_839, n_2_838, n_2_837, n_2_836, n_2_835, n_2_834, n_2_833, n_2_832, 
      n_2_831, n_2_778, n_2_777, n_2_776, n_2_775, n_2_774, n_2_773, n_2_772, 
      n_2_771, n_2_770, n_2_769, n_2_768, n_2_767, n_2_711, n_2_710, n_2_709, 
      n_2_708, n_2_707, n_2_706, n_2_705, n_2_704, n_2_703, n_2_9, n_2_8, n_2_7, 
      n_2_6, n_2_5, n_2_4, n_2_3, n_2_2, n_2_1, n_2_0, n_2_848, n_2_847, uc_817, 
      uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, uc_826, 
      uc_827, uc_828, uc_829, uc_830, uc_831, uc_832}), .carry_final());
   CSA__0_118 cs10 (.x({n_464, n_463, n_462, n_461, n_460, n_459, n_458, n_457, 
      n_456, n_455, n_454, n_453, n_452, n_451, n_450, n_449, n_448, n_447, 
      n_446, n_445, n_444, n_443, n_442, n_441, n_440, n_439, n_438, n_437, 
      n_436, n_435, n_434, n_433, n_432, n_431, n_430, n_429, n_428, n_427, 
      n_426, n_425, n_424, n_423, n_422, n_421, n_420, n_419, n_418, n_417, 
      n_416, n_415, n_414, n_413, n_412, n_411, n_410, n_409, n_408, n_407, 
      n_406, n_405, n_404, uc_833, uc_834, uc_835}), .y({n_524, n_523, n_522, 
      n_521, n_520, n_519, n_518, n_517, n_516, n_515, n_514, n_513, n_512, 
      n_511, n_510, n_509, n_508, n_507, n_506, n_505, n_504, n_503, n_502, 
      n_501, n_500, n_499, n_498, n_497, n_496, n_495, n_494, n_493, n_492, 
      n_491, n_490, n_489, n_488, n_487, n_486, n_485, n_484, n_483, n_482, 
      n_481, n_480, n_479, n_478, n_477, n_476, n_475, n_474, n_473, n_472, 
      n_471, n_470, n_469, n_468, n_467, n_466, n_465, n_161, uc_836, uc_837, 
      uc_838}), .z({n_581, n_580, n_579, n_578, n_577, n_576, n_575, n_574, 
      n_573, n_572, n_571, n_570, n_569, n_568, n_567, n_566, n_565, n_564, 
      n_563, n_562, n_561, n_560, n_559, n_558, n_557, n_556, n_555, n_554, 
      n_553, n_552, n_551, n_550, n_549, n_548, n_547, n_546, n_545, n_544, 
      n_543, n_542, n_541, n_540, n_539, n_538, n_537, n_536, n_535, n_534, 
      n_533, n_532, n_531, n_530, n_529, n_528, n_527, n_526, n_525, n_162, 
      uc_839, uc_840, uc_841, uc_842, uc_843, uc_844}), .s({n_694, n_693, n_692, 
      n_691, n_690, n_689, n_688, n_687, n_686, n_685, n_684, n_683, n_682, 
      n_681, n_680, n_679, n_678, n_677, n_676, n_675, n_674, n_673, n_672, 
      n_671, n_670, n_669, n_668, n_667, n_666, n_665, n_664, n_663, n_662, 
      n_661, n_660, n_659, n_658, n_657, n_656, n_655, n_654, n_653, n_652, 
      n_651, n_650, n_649, n_648, n_647, n_646, n_645, n_644, n_643, n_642, 
      n_641, n_640, n_639, n_638, n_637, n_636, n_635, n_634, uc_845, uc_846, 
      uc_847}), .carry_final());
   CSA__0_125 cs8 (.x({n_292, uc_848, uc_849, uc_850, uc_851, uc_852, uc_853, 
      uc_854, uc_855, n_291, n_290, n_289, n_288, n_287, n_286, n_285, n_284, 
      n_283, n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, 
      n_273, n_272, n_271, n_270, n_269, n_268, n_267, n_266, n_265, n_264, 
      n_263, n_262, uc_856, uc_857, uc_858, uc_859, uc_860, uc_861, uc_862, 
      uc_863, uc_864, uc_865, uc_866, uc_867, uc_868, uc_869, uc_870, uc_871, 
      uc_872, uc_873, uc_874, uc_875, uc_876, uc_877, uc_878, uc_879, uc_880}), 
      .y({n_324, uc_881, uc_882, uc_883, uc_884, uc_885, uc_886, uc_887, n_323, 
      n_322, n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314, n_313, 
      n_312, n_311, n_310, n_309, n_308, n_307, n_306, n_305, n_304, n_303, 
      n_302, n_301, n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, 
      uc_888, uc_889, uc_890, uc_891, uc_892, uc_893, uc_894, uc_895, uc_896, 
      uc_897, uc_898, uc_899, uc_900, uc_901, uc_902, uc_903, uc_904, uc_905, 
      uc_906, uc_907, uc_908, uc_909, uc_910, uc_911, uc_912}), .z({n_356, 
      uc_913, uc_914, uc_915, uc_916, uc_917, uc_918, n_355, n_354, n_353, n_352, 
      n_351, n_350, n_349, n_348, n_347, n_346, n_345, n_344, n_343, n_342, 
      n_341, n_340, n_339, n_338, n_337, n_336, n_335, n_334, n_333, n_332, 
      n_331, n_330, n_329, n_328, n_327, n_326, n_325, uc_919, uc_920, uc_921, 
      uc_922, uc_923, uc_924, uc_925, uc_926, uc_927, uc_928, uc_929, uc_930, 
      uc_931, uc_932, uc_933, uc_934, uc_935, uc_936, uc_937, uc_938, uc_939, 
      uc_940, uc_941, uc_942, uc_943, uc_944}), .s({n_733, n_732, n_731, n_730, 
      n_729, n_728, n_727, n_726, n_725, n_724, n_723, n_722, n_721, n_720, 
      n_719, n_718, n_717, n_716, n_715, n_714, n_713, n_712, n_711, n_710, 
      n_709, n_708, n_707, n_706, n_705, n_704, n_703, n_702, n_701, n_700, 
      n_699, n_698, n_697, n_696, n_695, uc_945, uc_946, uc_947, uc_948, uc_949, 
      uc_950, uc_951, uc_952, uc_953, uc_954, uc_955, uc_956, uc_957, uc_958, 
      uc_959, uc_960, uc_961, uc_962, uc_963, uc_964, uc_965, uc_966, uc_967, 
      uc_968, uc_969}), .carry_final());
   CSA__4_2043 cs7 (.x({n_196, uc_970, uc_971, uc_972, uc_973, uc_974, uc_975, 
      uc_976, uc_977, uc_978, uc_979, uc_980, n_195, n_194, n_193, n_192, n_191, 
      n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, 
      n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, 
      n_170, n_169, n_168, n_167, n_166, uc_981, uc_982, uc_983, uc_984, uc_985, 
      uc_986, uc_987, uc_988, uc_989, uc_990, uc_991, uc_992, uc_993, uc_994, 
      uc_995, uc_996, uc_997, uc_998, uc_999, uc_1000, uc_1001, uc_1002}), 
      .y({n_228, uc_1003, uc_1004, uc_1005, uc_1006, uc_1007, uc_1008, uc_1009, 
      uc_1010, uc_1011, uc_1012, n_227, n_226, n_225, n_224, n_223, n_222, n_221, 
      n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, 
      n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, n_201, 
      n_200, n_199, n_198, n_197, uc_1013, uc_1014, uc_1015, uc_1016, uc_1017, 
      uc_1018, uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, uc_1024, uc_1025, 
      uc_1026, uc_1027, uc_1028, uc_1029, uc_1030, uc_1031, uc_1032, uc_1033, 
      uc_1034}), .z({n_260, uc_1035, uc_1036, uc_1037, uc_1038, uc_1039, uc_1040, 
      uc_1041, uc_1042, uc_1043, n_259, n_258, n_257, n_256, n_255, n_254, n_253, 
      n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, 
      n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, 
      n_232, n_231, n_230, n_229, uc_1044, uc_1045, uc_1046, uc_1047, uc_1048, 
      uc_1049, uc_1050, uc_1051, uc_1052, uc_1053, uc_1054, uc_1055, uc_1056, 
      uc_1057, uc_1058, uc_1059, uc_1060, uc_1061, uc_1062, uc_1063, uc_1064, 
      uc_1065, uc_1066}), .s({n_5_63, n_5_62, n_5_61, n_5_60, n_5_59, n_5_58, 
      n_5_57, n_5_56, n_5_55, n_5_54, n_5_53, n_5_52, n_5_51, n_5_50, n_5_49, 
      n_5_48, n_5_47, n_5_46, n_5_45, n_5_44, n_5_43, n_5_42, n_5_41, n_5_40, 
      n_5_39, n_5_38, n_5_37, n_5_36, n_5_35, n_5_34, n_5_33, n_5_32, n_5_31, 
      n_5_30, n_5_29, n_5_28, n_5_27, n_5_26, n_5_25, n_5_24, n_5_23, n_5_22, 
      uc_1067, uc_1068, uc_1069, uc_1070, uc_1071, uc_1072, uc_1073, uc_1074, 
      uc_1075, uc_1076, uc_1077, uc_1078, uc_1079, uc_1080, uc_1081, uc_1082, 
      uc_1083, uc_1084, uc_1085, uc_1086, uc_1087, uc_1088}), .carry_final());
   CSA__4_3068 cs14 (.x({n_694, n_693, n_692, n_691, n_690, n_689, n_688, n_687, 
      n_686, n_685, n_684, n_683, n_682, n_681, n_680, n_679, n_678, n_677, 
      n_676, n_675, n_674, n_673, n_672, n_671, n_670, n_669, n_668, n_667, 
      n_666, n_665, n_664, n_663, n_662, n_661, n_660, n_659, n_658, n_657, 
      n_656, n_655, n_654, n_653, n_652, n_651, n_650, n_649, n_648, n_647, 
      n_646, n_645, n_644, n_643, n_642, n_641, n_640, uc_1089, uc_1090, uc_1091, 
      uc_1092, uc_1093, uc_1094, uc_1095, uc_1096, uc_1097}), .y({n_633, n_632, 
      n_631, n_630, n_629, n_628, n_627, n_626, n_625, n_624, n_623, n_622, 
      n_621, n_620, n_619, n_618, n_617, n_616, n_615, n_614, n_613, n_612, 
      n_611, n_610, n_609, n_608, n_607, n_606, n_605, n_604, n_603, n_602, 
      n_601, n_600, n_599, n_598, n_597, n_596, n_595, n_594, n_593, n_592, 
      n_591, n_590, n_589, n_588, n_587, n_586, n_585, n_584, n_583, n_582, 
      n_2_714__1, n_2_713__1, n_163, uc_1098, uc_1099, uc_1100, uc_1101, uc_1102, 
      uc_1103, uc_1104, uc_1105, uc_1106}), .z({n_5_84, n_5_83, n_5_82, n_5_81, 
      n_5_80, n_5_79, n_5_78, n_5_77, n_5_76, n_5_75, n_5_74, n_5_73, n_5_72, 
      n_5_71, n_5_70, n_5_69, n_5_68, n_5_67, n_5_66, n_5_65, n_5_64, n_5_21, 
      n_5_20, n_5_19, n_5_18, n_5_17, n_5_16, n_5_15, n_5_14, n_5_13, n_5_12, 
      n_5_11, n_5_10, n_5_9, n_5_8, n_5_7, n_5_6, n_5_5, n_5_4, n_5_3, n_5_2, 
      n_5_1, n_5_0, n_358, n_357, n_164, uc_1107, uc_1108, uc_1109, uc_1110, 
      uc_1111, uc_1112, uc_1113, uc_1114, uc_1115, uc_1116, uc_1117, uc_1118, 
      uc_1119, uc_1120, uc_1121, uc_1122, uc_1123, uc_1124}), .s({n_788, n_787, 
      n_786, n_785, n_784, n_783, n_782, n_781, n_780, n_779, n_778, n_777, 
      n_776, n_775, n_774, n_773, n_772, n_771, n_770, n_769, n_768, n_767, 
      n_766, n_765, n_764, n_763, n_762, n_761, n_760, n_759, n_758, n_757, 
      n_756, n_755, n_754, n_753, n_752, n_751, n_750, n_749, n_748, n_747, 
      n_746, n_745, n_744, n_743, n_742, n_741, n_740, n_739, n_738, n_737, 
      n_736, n_735, n_734, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, uc_1130, 
      uc_1131, uc_1132, uc_1133}), .carry_final());
   CSA__0_131 cs12 (.x({n_401, n_400, n_399, n_398, n_397, n_396, n_395, n_394, 
      n_393, n_392, n_391, n_390, n_389, n_388, n_387, n_386, n_385, n_384, 
      n_383, n_382, n_381, n_380, n_379, n_378, n_377, n_376, n_375, n_374, 
      n_373, n_372, n_371, n_370, n_369, n_368, n_367, n_366, n_365, n_364, 
      n_363, n_362, n_361, n_360, n_359, uc_1134, uc_1135, uc_1136, uc_1137, 
      uc_1138, uc_1139, uc_1140, uc_1141, uc_1142, uc_1143, uc_1144, uc_1145, 
      uc_1146, uc_1147, uc_1148, uc_1149, uc_1150, uc_1151, uc_1152, uc_1153, 
      uc_1154}), .y({n_5_63, n_5_62, n_5_61, n_5_60, n_5_59, n_5_58, n_5_57, 
      n_5_56, n_5_55, n_5_54, n_5_53, n_5_52, n_5_51, n_5_50, n_5_49, n_5_48, 
      n_5_47, n_5_46, n_5_45, n_5_44, n_5_43, n_5_42, n_5_41, n_5_40, n_5_39, 
      n_5_38, n_5_37, n_5_36, n_5_35, n_5_34, n_5_33, n_5_32, n_5_31, n_5_30, 
      n_5_29, n_5_28, n_5_27, n_5_26, n_5_25, n_5_24, n_5_23, n_5_22, n_165, 
      uc_1155, uc_1156, uc_1157, uc_1158, uc_1159, uc_1160, uc_1161, uc_1162, 
      uc_1163, uc_1164, uc_1165, uc_1166, uc_1167, uc_1168, uc_1169, uc_1170, 
      uc_1171, uc_1172, uc_1173, uc_1174, uc_1175}), .z({n_733, n_732, n_731, 
      n_730, n_729, n_728, n_727, n_726, n_725, n_724, n_723, n_722, n_721, 
      n_720, n_719, n_718, n_717, n_716, n_715, n_714, n_713, n_712, n_711, 
      n_710, n_709, n_708, n_707, n_706, n_705, n_704, n_703, n_702, n_701, 
      n_700, n_699, n_698, n_697, n_696, n_695, n_261, uc_1176, uc_1177, uc_1178, 
      uc_1179, uc_1180, uc_1181, uc_1182, uc_1183, uc_1184, uc_1185, uc_1186, 
      uc_1187, uc_1188, uc_1189, uc_1190, uc_1191, uc_1192, uc_1193, uc_1194, 
      uc_1195, uc_1196, uc_1197, uc_1198, uc_1199}), .s({n_5_84, n_5_83, n_5_82, 
      n_5_81, n_5_80, n_5_79, n_5_78, n_5_77, n_5_76, n_5_75, n_5_74, n_5_73, 
      n_5_72, n_5_71, n_5_70, n_5_69, n_5_68, n_5_67, n_5_66, n_5_65, n_5_64, 
      n_5_21, n_5_20, n_5_19, n_5_18, n_5_17, n_5_16, n_5_15, n_5_14, n_5_13, 
      n_5_12, n_5_11, n_5_10, n_5_9, n_5_8, n_5_7, n_5_6, n_5_5, n_5_4, n_5_3, 
      n_5_2, n_5_1, n_5_0, uc_1200, uc_1201, uc_1202, uc_1203, uc_1204, uc_1205, 
      uc_1206, uc_1207, uc_1208, uc_1209, uc_1210, uc_1211, uc_1212, uc_1213, 
      uc_1214, uc_1215, uc_1216, uc_1217, uc_1218, uc_1219, uc_1220}), 
      .carry_final());
   CSA__5_2043 cs13 (.x({n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, 
      n_0_93, n_0_92, n_0_91, n_0_64, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, 
      n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, 
      n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, 
      n_0_67, uc_1221, uc_1222, uc_1223, uc_1224, uc_1225, uc_1226, uc_1227, 
      uc_1228, uc_1229, uc_1230, uc_1231, uc_1232, uc_1233, uc_1234, uc_1235, 
      uc_1236, uc_1237, uc_1238, uc_1239, uc_1240, uc_1241, uc_1242, uc_1243, 
      uc_1244, uc_1245, uc_1246, uc_1247, uc_1248, uc_1249, uc_1250}), .y({n_127, 
      uc_1251, uc_1252, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, 
      n_118, n_117, n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, 
      n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
      n_97, n_96, uc_1253, uc_1254, uc_1255, uc_1256, uc_1257, uc_1258, uc_1259, 
      uc_1260, uc_1261, uc_1262, uc_1263, uc_1264, uc_1265, uc_1266, uc_1267, 
      uc_1268, uc_1269, uc_1270, uc_1271, uc_1272, uc_1273, uc_1274, uc_1275, 
      uc_1276, uc_1277, uc_1278, uc_1279, uc_1280, uc_1281, uc_1282}), .z({n_159, 
      uc_1283, n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, n_150, 
      n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, n_140, 
      n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, n_130, 
      n_129, n_128, uc_1284, uc_1285, uc_1286, uc_1287, uc_1288, uc_1289, 
      uc_1290, uc_1291, uc_1292, uc_1293, uc_1294, uc_1295, uc_1296, uc_1297, 
      uc_1298, uc_1299, uc_1300, uc_1301, uc_1302, uc_1303, uc_1304, uc_1305, 
      uc_1306, uc_1307, uc_1308, uc_1309, uc_1310, uc_1311, uc_1312, uc_1313, 
      uc_1314}), .s({n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, 
      n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, 
      n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, 
      n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, 
      n_0_97, n_0_96, n_0_95, n_0_94, uc_1315, uc_1316, uc_1317, uc_1318, 
      uc_1319, uc_1320, uc_1321, uc_1322, uc_1323, uc_1324, uc_1325, uc_1326, 
      uc_1327, uc_1328, uc_1329, uc_1330, uc_1331, uc_1332, uc_1333, uc_1334, 
      uc_1335, uc_1336, uc_1337, uc_1338, uc_1339, uc_1340, uc_1341, uc_1342, 
      uc_1343, uc_1344}), .carry_final());
   carry_increment_adder ci (.in1({n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, 
      n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, 
      n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, 
      n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, 
      n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_66, n_0_65, n_0, uc_1345, 
      uc_1346, uc_1347, uc_1348, uc_1349, uc_1350, uc_1351, uc_1352, uc_1353, 
      uc_1354, uc_1355, uc_1356, uc_1357, uc_1358, uc_1359, uc_1360, uc_1361, 
      uc_1362, uc_1363, uc_1364, uc_1365, uc_1366, uc_1367, uc_1368, uc_1369, 
      uc_1370, uc_1371}), .in2({n_788, n_787, n_786, n_785, n_784, n_783, n_782, 
      n_781, n_780, n_779, n_778, n_777, n_776, n_775, n_774, n_773, n_772, 
      n_771, n_770, n_769, n_768, n_767, n_766, n_765, n_764, n_763, n_762, 
      n_761, n_760, n_759, n_758, n_757, n_756, n_755, n_754, n_753, n_752, 
      uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, uc_1377, uc_1378, uc_1379, 
      uc_1380, uc_1381, uc_1382, uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, 
      uc_1388, uc_1389, uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, 
      uc_1396, uc_1397, uc_1398}), .s({product[63], product[62], product[61], 
      product[60], product[59], product[58], product[57], product[56], 
      product[55], product[54], product[53], product[52], product[51], 
      product[50], product[49], product[48], product[47], product[46], 
      product[45], product[44], product[43], product[42], product[41], 
      product[40], product[39], product[38], product[37], product[36], 
      product[35], product[34], product[33], product[32], product[31], 
      product[30], product[29], product[28], product[27], uc_1399, uc_1400, 
      uc_1401, uc_1402, uc_1403, uc_1404, uc_1405, uc_1406, uc_1407, uc_1408, 
      uc_1409, uc_1410, uc_1411, uc_1412, uc_1413, uc_1414, uc_1415, uc_1416, 
      uc_1417, uc_1418, uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, uc_1424, 
      uc_1425}), .cin(), .cout(), .OF());
   DFF_X1 \Out_reg[63]  (.D(n_0_128), .CK(clk), .Q(Out[63]), .QN());
   DFF_X1 \Out_reg[62]  (.D(n_0_63), .CK(clk), .Q(Out[62]), .QN());
   DFF_X1 \Out_reg[61]  (.D(n_0_62), .CK(clk), .Q(Out[61]), .QN());
   DFF_X1 \Out_reg[60]  (.D(n_0_61), .CK(clk), .Q(Out[60]), .QN());
   DFF_X1 \Out_reg[59]  (.D(n_0_60), .CK(clk), .Q(Out[59]), .QN());
   DFF_X1 \Out_reg[58]  (.D(n_0_59), .CK(clk), .Q(Out[58]), .QN());
   DFF_X1 \Out_reg[57]  (.D(n_0_58), .CK(clk), .Q(Out[57]), .QN());
   DFF_X1 \Out_reg[56]  (.D(n_0_57), .CK(clk), .Q(Out[56]), .QN());
   DFF_X1 \Out_reg[55]  (.D(n_0_56), .CK(clk), .Q(Out[55]), .QN());
   DFF_X1 \Out_reg[54]  (.D(n_0_55), .CK(clk), .Q(Out[54]), .QN());
   DFF_X1 \Out_reg[53]  (.D(n_0_54), .CK(clk), .Q(Out[53]), .QN());
   DFF_X1 \Out_reg[52]  (.D(n_0_53), .CK(clk), .Q(Out[52]), .QN());
   DFF_X1 \Out_reg[51]  (.D(n_0_52), .CK(clk), .Q(Out[51]), .QN());
   DFF_X1 \Out_reg[50]  (.D(n_0_51), .CK(clk), .Q(Out[50]), .QN());
   DFF_X1 \Out_reg[49]  (.D(n_0_50), .CK(clk), .Q(Out[49]), .QN());
   DFF_X1 \Out_reg[48]  (.D(n_0_49), .CK(clk), .Q(Out[48]), .QN());
   DFF_X1 \Out_reg[47]  (.D(n_0_48), .CK(clk), .Q(Out[47]), .QN());
   DFF_X1 \Out_reg[46]  (.D(n_0_47), .CK(clk), .Q(Out[46]), .QN());
   DFF_X1 \Out_reg[45]  (.D(n_0_46), .CK(clk), .Q(Out[45]), .QN());
   DFF_X1 \Out_reg[44]  (.D(n_0_45), .CK(clk), .Q(Out[44]), .QN());
   DFF_X1 \Out_reg[43]  (.D(n_0_44), .CK(clk), .Q(Out[43]), .QN());
   DFF_X1 \Out_reg[42]  (.D(n_0_43), .CK(clk), .Q(Out[42]), .QN());
   DFF_X1 \Out_reg[41]  (.D(n_0_42), .CK(clk), .Q(Out[41]), .QN());
   DFF_X1 \Out_reg[40]  (.D(n_0_41), .CK(clk), .Q(Out[40]), .QN());
   DFF_X1 \Out_reg[39]  (.D(n_0_40), .CK(clk), .Q(Out[39]), .QN());
   DFF_X1 \Out_reg[38]  (.D(n_0_39), .CK(clk), .Q(Out[38]), .QN());
   DFF_X1 \Out_reg[37]  (.D(n_0_38), .CK(clk), .Q(Out[37]), .QN());
   DFF_X1 \Out_reg[36]  (.D(n_0_37), .CK(clk), .Q(Out[36]), .QN());
   DFF_X1 \Out_reg[35]  (.D(n_0_36), .CK(clk), .Q(Out[35]), .QN());
   DFF_X1 \Out_reg[34]  (.D(n_0_35), .CK(clk), .Q(Out[34]), .QN());
   DFF_X1 \Out_reg[33]  (.D(n_0_34), .CK(clk), .Q(Out[33]), .QN());
   DFF_X1 \Out_reg[32]  (.D(n_0_33), .CK(clk), .Q(Out[32]), .QN());
   DFF_X1 \Out_reg[31]  (.D(n_0_32), .CK(clk), .Q(Out[31]), .QN());
   DFF_X1 \Out_reg[30]  (.D(n_0_31), .CK(clk), .Q(Out[30]), .QN());
   DFF_X1 \Out_reg[29]  (.D(n_0_30), .CK(clk), .Q(Out[29]), .QN());
   DFF_X1 \Out_reg[28]  (.D(n_0_29), .CK(clk), .Q(Out[28]), .QN());
   DFF_X1 \Out_reg[27]  (.D(n_0_28), .CK(clk), .Q(Out[27]), .QN());
   DFF_X1 \Out_reg[26]  (.D(n_0_27), .CK(clk), .Q(Out[26]), .QN());
   DFF_X1 \Out_reg[25]  (.D(n_0_26), .CK(clk), .Q(Out[25]), .QN());
   DFF_X1 \Out_reg[24]  (.D(n_0_25), .CK(clk), .Q(Out[24]), .QN());
   DFF_X1 \Out_reg[23]  (.D(n_0_24), .CK(clk), .Q(Out[23]), .QN());
   DFF_X1 \Out_reg[22]  (.D(n_0_23), .CK(clk), .Q(Out[22]), .QN());
   DFF_X1 \Out_reg[21]  (.D(n_0_22), .CK(clk), .Q(Out[21]), .QN());
   DFF_X1 \Out_reg[20]  (.D(n_0_21), .CK(clk), .Q(Out[20]), .QN());
   DFF_X1 \Out_reg[19]  (.D(n_0_20), .CK(clk), .Q(Out[19]), .QN());
   DFF_X1 \Out_reg[18]  (.D(n_0_19), .CK(clk), .Q(Out[18]), .QN());
   DFF_X1 \Out_reg[17]  (.D(n_0_18), .CK(clk), .Q(Out[17]), .QN());
   DFF_X1 \Out_reg[16]  (.D(n_0_17), .CK(clk), .Q(Out[16]), .QN());
   DFF_X1 \Out_reg[15]  (.D(n_0_16), .CK(clk), .Q(Out[15]), .QN());
   DFF_X1 \Out_reg[14]  (.D(n_0_15), .CK(clk), .Q(Out[14]), .QN());
   DFF_X1 \Out_reg[13]  (.D(n_0_14), .CK(clk), .Q(Out[13]), .QN());
   DFF_X1 \Out_reg[12]  (.D(n_0_13), .CK(clk), .Q(Out[12]), .QN());
   DFF_X1 \Out_reg[11]  (.D(n_0_12), .CK(clk), .Q(Out[11]), .QN());
   DFF_X1 \Out_reg[10]  (.D(n_0_11), .CK(clk), .Q(Out[10]), .QN());
   DFF_X1 \Out_reg[9]  (.D(n_0_10), .CK(clk), .Q(Out[9]), .QN());
   DFF_X1 \Out_reg[8]  (.D(n_0_9), .CK(clk), .Q(Out[8]), .QN());
   DFF_X1 \Out_reg[7]  (.D(n_0_8), .CK(clk), .Q(Out[7]), .QN());
   DFF_X1 \Out_reg[6]  (.D(n_0_7), .CK(clk), .Q(Out[6]), .QN());
   DFF_X1 \Out_reg[5]  (.D(n_0_6), .CK(clk), .Q(Out[5]), .QN());
   DFF_X1 \Out_reg[4]  (.D(n_0_5), .CK(clk), .Q(Out[4]), .QN());
   DFF_X1 \Out_reg[3]  (.D(n_0_4), .CK(clk), .Q(Out[3]), .QN());
   DFF_X1 \Out_reg[2]  (.D(n_0_3), .CK(clk), .Q(Out[2]), .QN());
   DFF_X1 \Out_reg[1]  (.D(n_0_2), .CK(clk), .Q(Out[1]), .QN());
   DFF_X1 \Out_reg[0]  (.D(n_0_1), .CK(clk), .Q(Out[0]), .QN());
   DFF_X1 \y_reg[26]  (.D(B[26]), .CK(n_0_129), .Q(y), .QN());
   DFF_X1 \y_reg[25]  (.D(B[25]), .CK(n_0_129), .Q(n_789), .QN());
   DFF_X1 \y_reg[24]  (.D(B[24]), .CK(n_0_129), .Q(n_790), .QN());
   DFF_X1 \y_reg[23]  (.D(B[23]), .CK(n_0_129), .Q(n_791), .QN());
   DFF_X1 \y_reg[22]  (.D(B[22]), .CK(n_0_129), .Q(n_792), .QN());
   DFF_X1 \y_reg[21]  (.D(B[21]), .CK(n_0_129), .Q(n_793), .QN());
   DFF_X1 \y_reg[20]  (.D(B[20]), .CK(n_0_129), .Q(n_794), .QN());
   DFF_X1 \y_reg[19]  (.D(B[19]), .CK(n_0_129), .Q(n_795), .QN());
   DFF_X1 \y_reg[18]  (.D(B[18]), .CK(n_0_129), .Q(n_796), .QN());
   DFF_X1 \y_reg[17]  (.D(B[17]), .CK(n_0_129), .Q(n_797), .QN());
   DFF_X1 \y_reg[16]  (.D(B[16]), .CK(n_0_129), .Q(n_798), .QN());
   DFF_X1 \y_reg[15]  (.D(B[15]), .CK(n_0_129), .Q(n_799), .QN());
   DFF_X1 \y_reg[14]  (.D(B[14]), .CK(n_0_129), .Q(n_800), .QN());
   DFF_X1 \y_reg[13]  (.D(B[13]), .CK(n_0_129), .Q(n_801), .QN());
   DFF_X1 \y_reg[12]  (.D(B[12]), .CK(n_0_129), .Q(n_802), .QN());
   DFF_X1 \y_reg[11]  (.D(B[11]), .CK(n_0_129), .Q(n_803), .QN());
   DFF_X1 \y_reg[10]  (.D(B[10]), .CK(n_0_129), .Q(n_804), .QN());
   DFF_X1 \y_reg[9]  (.D(B[9]), .CK(n_0_129), .Q(n_805), .QN());
   DFF_X1 \y_reg[8]  (.D(B[8]), .CK(n_0_129), .Q(n_806), .QN());
   DFF_X1 \y_reg[7]  (.D(B[7]), .CK(n_0_129), .Q(n_807), .QN());
   DFF_X1 \y_reg[6]  (.D(B[6]), .CK(n_0_129), .Q(n_808), .QN());
   DFF_X1 \y_reg[5]  (.D(B[5]), .CK(n_0_129), .Q(n_809), .QN());
   DFF_X1 \y_reg[4]  (.D(B[4]), .CK(n_0_129), .Q(n_810), .QN());
   DFF_X1 \y_reg[3]  (.D(B[3]), .CK(n_0_129), .Q(n_811), .QN());
   DFF_X1 \y_reg[2]  (.D(B[2]), .CK(n_0_129), .Q(n_812), .QN());
   DFF_X1 \y_reg[1]  (.D(B[1]), .CK(n_0_129), .Q(n_813), .QN());
   DFF_X1 \y_reg[0]  (.D(B[0]), .CK(n_0_129), .Q(n_814), .QN());
   DFF_X1 \y_reg[31]  (.D(B[31]), .CK(n_0_129), .Q(n_815), .QN());
   DFF_X1 \y_reg[30]  (.D(B[30]), .CK(n_0_129), .Q(n_816), .QN());
   DFF_X1 \y_reg[29]  (.D(B[29]), .CK(n_0_129), .Q(n_817), .QN());
   DFF_X1 \y_reg[28]  (.D(B[28]), .CK(n_0_129), .Q(n_818), .QN());
   DFF_X1 \x_reg[31]  (.D(A[31]), .CK(n_0_129), .Q(x[31]), .QN());
   DFF_X1 \x_reg[30]  (.D(A[30]), .CK(n_0_129), .Q(x[30]), .QN());
   DFF_X1 \x_reg[29]  (.D(A[29]), .CK(n_0_129), .Q(x[29]), .QN());
   DFF_X1 \x_reg[28]  (.D(A[28]), .CK(n_0_129), .Q(x[28]), .QN());
   DFF_X1 \x_reg[27]  (.D(A[27]), .CK(n_0_129), .Q(x[27]), .QN());
   DFF_X1 \x_reg[26]  (.D(A[26]), .CK(n_0_129), .Q(x[26]), .QN());
   DFF_X1 \x_reg[25]  (.D(A[25]), .CK(n_0_129), .Q(x[25]), .QN());
   DFF_X1 \x_reg[24]  (.D(A[24]), .CK(n_0_129), .Q(x[24]), .QN());
   DFF_X1 \x_reg[23]  (.D(A[23]), .CK(n_0_129), .Q(x[23]), .QN());
   DFF_X1 \x_reg[22]  (.D(A[22]), .CK(n_0_129), .Q(x[22]), .QN());
   DFF_X1 \x_reg[21]  (.D(A[21]), .CK(n_0_129), .Q(x[21]), .QN());
   DFF_X1 \x_reg[20]  (.D(A[20]), .CK(n_0_129), .Q(x[20]), .QN());
   DFF_X1 \x_reg[19]  (.D(A[19]), .CK(n_0_129), .Q(x[19]), .QN());
   DFF_X1 \x_reg[18]  (.D(A[18]), .CK(n_0_129), .Q(x[18]), .QN());
   DFF_X1 \x_reg[17]  (.D(A[17]), .CK(n_0_129), .Q(x[17]), .QN());
   DFF_X1 \x_reg[16]  (.D(A[16]), .CK(n_0_129), .Q(x[16]), .QN());
   DFF_X1 \x_reg[15]  (.D(A[15]), .CK(n_0_129), .Q(x[15]), .QN());
   DFF_X1 \x_reg[14]  (.D(A[14]), .CK(n_0_129), .Q(x[14]), .QN());
   DFF_X1 \x_reg[13]  (.D(A[13]), .CK(n_0_129), .Q(x[13]), .QN());
   DFF_X1 \x_reg[12]  (.D(A[12]), .CK(n_0_129), .Q(x[12]), .QN());
   DFF_X1 \x_reg[11]  (.D(A[11]), .CK(n_0_129), .Q(x[11]), .QN());
   DFF_X1 \x_reg[10]  (.D(A[10]), .CK(n_0_129), .Q(x[10]), .QN());
   DFF_X1 \x_reg[9]  (.D(A[9]), .CK(n_0_129), .Q(x[9]), .QN());
   DFF_X1 \x_reg[8]  (.D(A[8]), .CK(n_0_129), .Q(x[8]), .QN());
   DFF_X1 \x_reg[7]  (.D(A[7]), .CK(n_0_129), .Q(x[7]), .QN());
   DFF_X1 \x_reg[6]  (.D(A[6]), .CK(n_0_129), .Q(x[6]), .QN());
   DFF_X1 \x_reg[5]  (.D(A[5]), .CK(n_0_129), .Q(x[5]), .QN());
   DFF_X1 \x_reg[4]  (.D(A[4]), .CK(n_0_129), .Q(x[4]), .QN());
   DFF_X1 \x_reg[3]  (.D(A[3]), .CK(n_0_129), .Q(x[3]), .QN());
   DFF_X1 \x_reg[2]  (.D(A[2]), .CK(n_0_129), .Q(x[2]), .QN());
   DFF_X1 \x_reg[1]  (.D(A[1]), .CK(n_0_129), .Q(x[1]), .QN());
   DFF_X1 \x_reg[0]  (.D(A[0]), .CK(n_0_129), .Q(x[0]), .QN());
   DFF_X1 \y_reg[27]  (.D(B[27]), .CK(n_0_129), .Q(n_819), .QN());
   INV_X1 i_0_0_0 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_0_1 (.A1(n_0_0), .A2(n_160), .ZN(n_0_1));
   AND2_X1 i_0_0_2 (.A1(n_0_0), .A2(n_402), .ZN(n_0_2));
   AND2_X1 i_0_0_3 (.A1(n_0_0), .A2(n_403), .ZN(n_0_3));
   AND2_X1 i_0_0_4 (.A1(n_0_0), .A2(n_634), .ZN(n_0_4));
   AND2_X1 i_0_0_5 (.A1(n_0_0), .A2(n_635), .ZN(n_0_5));
   AND2_X1 i_0_0_6 (.A1(n_0_0), .A2(n_636), .ZN(n_0_6));
   AND2_X1 i_0_0_7 (.A1(n_0_0), .A2(n_637), .ZN(n_0_7));
   AND2_X1 i_0_0_8 (.A1(n_0_0), .A2(n_638), .ZN(n_0_8));
   AND2_X1 i_0_0_9 (.A1(n_0_0), .A2(n_639), .ZN(n_0_9));
   AND2_X1 i_0_0_10 (.A1(n_0_0), .A2(n_734), .ZN(n_0_10));
   AND2_X1 i_0_0_11 (.A1(n_0_0), .A2(n_735), .ZN(n_0_11));
   AND2_X1 i_0_0_12 (.A1(n_0_0), .A2(n_736), .ZN(n_0_12));
   AND2_X1 i_0_0_13 (.A1(n_0_0), .A2(n_737), .ZN(n_0_13));
   AND2_X1 i_0_0_14 (.A1(n_0_0), .A2(n_738), .ZN(n_0_14));
   AND2_X1 i_0_0_15 (.A1(n_0_0), .A2(n_739), .ZN(n_0_15));
   AND2_X1 i_0_0_16 (.A1(n_0_0), .A2(n_740), .ZN(n_0_16));
   AND2_X1 i_0_0_17 (.A1(n_0_0), .A2(n_741), .ZN(n_0_17));
   AND2_X1 i_0_0_18 (.A1(n_0_0), .A2(n_742), .ZN(n_0_18));
   AND2_X1 i_0_0_19 (.A1(n_0_0), .A2(n_743), .ZN(n_0_19));
   AND2_X1 i_0_0_20 (.A1(n_0_0), .A2(n_744), .ZN(n_0_20));
   AND2_X1 i_0_0_21 (.A1(n_0_0), .A2(n_745), .ZN(n_0_21));
   AND2_X1 i_0_0_22 (.A1(n_0_0), .A2(n_746), .ZN(n_0_22));
   AND2_X1 i_0_0_23 (.A1(n_0_0), .A2(n_747), .ZN(n_0_23));
   AND2_X1 i_0_0_24 (.A1(n_0_0), .A2(n_748), .ZN(n_0_24));
   AND2_X1 i_0_0_25 (.A1(n_0_0), .A2(n_749), .ZN(n_0_25));
   AND2_X1 i_0_0_26 (.A1(n_0_0), .A2(n_750), .ZN(n_0_26));
   AND2_X1 i_0_0_27 (.A1(n_0_0), .A2(n_751), .ZN(n_0_27));
   AND2_X1 i_0_0_28 (.A1(n_0_0), .A2(product[27]), .ZN(n_0_28));
   AND2_X1 i_0_0_29 (.A1(n_0_0), .A2(product[28]), .ZN(n_0_29));
   AND2_X1 i_0_0_30 (.A1(n_0_0), .A2(product[29]), .ZN(n_0_30));
   AND2_X1 i_0_0_31 (.A1(n_0_0), .A2(product[30]), .ZN(n_0_31));
   AND2_X1 i_0_0_32 (.A1(n_0_0), .A2(product[31]), .ZN(n_0_32));
   AND2_X1 i_0_0_33 (.A1(n_0_0), .A2(product[32]), .ZN(n_0_33));
   AND2_X1 i_0_0_34 (.A1(n_0_0), .A2(product[33]), .ZN(n_0_34));
   AND2_X1 i_0_0_35 (.A1(n_0_0), .A2(product[34]), .ZN(n_0_35));
   AND2_X1 i_0_0_36 (.A1(n_0_0), .A2(product[35]), .ZN(n_0_36));
   AND2_X1 i_0_0_37 (.A1(n_0_0), .A2(product[36]), .ZN(n_0_37));
   AND2_X1 i_0_0_38 (.A1(n_0_0), .A2(product[37]), .ZN(n_0_38));
   AND2_X1 i_0_0_39 (.A1(n_0_0), .A2(product[38]), .ZN(n_0_39));
   AND2_X1 i_0_0_40 (.A1(n_0_0), .A2(product[39]), .ZN(n_0_40));
   AND2_X1 i_0_0_41 (.A1(n_0_0), .A2(product[40]), .ZN(n_0_41));
   AND2_X1 i_0_0_42 (.A1(n_0_0), .A2(product[41]), .ZN(n_0_42));
   AND2_X1 i_0_0_43 (.A1(n_0_0), .A2(product[42]), .ZN(n_0_43));
   AND2_X1 i_0_0_44 (.A1(n_0_0), .A2(product[43]), .ZN(n_0_44));
   AND2_X1 i_0_0_45 (.A1(n_0_0), .A2(product[44]), .ZN(n_0_45));
   AND2_X1 i_0_0_46 (.A1(n_0_0), .A2(product[45]), .ZN(n_0_46));
   AND2_X1 i_0_0_47 (.A1(n_0_0), .A2(product[46]), .ZN(n_0_47));
   AND2_X1 i_0_0_48 (.A1(n_0_0), .A2(product[47]), .ZN(n_0_48));
   AND2_X1 i_0_0_49 (.A1(n_0_0), .A2(product[48]), .ZN(n_0_49));
   AND2_X1 i_0_0_50 (.A1(n_0_0), .A2(product[49]), .ZN(n_0_50));
   AND2_X1 i_0_0_51 (.A1(n_0_0), .A2(product[50]), .ZN(n_0_51));
   AND2_X1 i_0_0_52 (.A1(n_0_0), .A2(product[51]), .ZN(n_0_52));
   AND2_X1 i_0_0_53 (.A1(n_0_0), .A2(product[52]), .ZN(n_0_53));
   AND2_X1 i_0_0_54 (.A1(n_0_0), .A2(product[53]), .ZN(n_0_54));
   AND2_X1 i_0_0_55 (.A1(n_0_0), .A2(product[54]), .ZN(n_0_55));
   AND2_X1 i_0_0_56 (.A1(n_0_0), .A2(product[55]), .ZN(n_0_56));
   AND2_X1 i_0_0_57 (.A1(n_0_0), .A2(product[56]), .ZN(n_0_57));
   AND2_X1 i_0_0_58 (.A1(n_0_0), .A2(product[57]), .ZN(n_0_58));
   AND2_X1 i_0_0_59 (.A1(n_0_0), .A2(product[58]), .ZN(n_0_59));
   AND2_X1 i_0_0_60 (.A1(n_0_0), .A2(product[59]), .ZN(n_0_60));
   AND2_X1 i_0_0_61 (.A1(n_0_0), .A2(product[60]), .ZN(n_0_61));
   AND2_X1 i_0_0_62 (.A1(n_0_0), .A2(product[61]), .ZN(n_0_62));
   AND2_X1 i_0_0_63 (.A1(n_0_0), .A2(product[62]), .ZN(n_0_63));
   AND2_X1 i_0_0_64 (.A1(n_0_0), .A2(product[63]), .ZN(n_0_128));
   CLKGATETST_X1 clk_gate_y_reg (.CK(clk), .E(n_0_0), .SE(1'b0), .GCK(n_0_129));
   CSA cs9 (.x({n_31, uc_1426, uc_1427, uc_1428, uc_1429, uc_1430, n_30, n_29, 
      n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
      n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, 
      n_3, n_2, n_1, uc_1431, uc_1432, uc_1433, uc_1434, uc_1435, uc_1436, 
      uc_1437, uc_1438, uc_1439, uc_1440, uc_1441, uc_1442, uc_1443, uc_1444, 
      uc_1445, uc_1446, uc_1447, uc_1448, uc_1449, uc_1450, uc_1451, uc_1452, 
      uc_1453, uc_1454, uc_1455, uc_1456, uc_1457, uc_1458}), .y({n_63, uc_1459, 
      uc_1460, uc_1461, uc_1462, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, 
      n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
      n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, uc_1463, 
      uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, uc_1469, uc_1470, uc_1471, 
      uc_1472, uc_1473, uc_1474, uc_1475, uc_1476, uc_1477, uc_1478, uc_1479, 
      uc_1480, uc_1481, uc_1482, uc_1483, uc_1484, uc_1485, uc_1486, uc_1487, 
      uc_1488, uc_1489, uc_1490}), .z({n_95, uc_1491, uc_1492, uc_1493, n_94, 
      n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, 
      n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, 
      n_69, n_68, n_67, n_66, n_65, n_64, uc_1494, uc_1495, uc_1496, uc_1497, 
      uc_1498, uc_1499, uc_1500, uc_1501, uc_1502, uc_1503, uc_1504, uc_1505, 
      uc_1506, uc_1507, uc_1508, uc_1509, uc_1510, uc_1511, uc_1512, uc_1513, 
      uc_1514, uc_1515, uc_1516, uc_1517, uc_1518, uc_1519, uc_1520, uc_1521, 
      uc_1522}), .s({n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, 
      n_0_93, n_0_92, n_0_91, n_0_64, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, 
      n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, 
      n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, 
      n_0_67, n_0_66, n_0_65, uc_1523, uc_1524, uc_1525, uc_1526, uc_1527, 
      uc_1528, uc_1529, uc_1530, uc_1531, uc_1532, uc_1533, uc_1534, uc_1535, 
      uc_1536, uc_1537, uc_1538, uc_1539, uc_1540, uc_1541, uc_1542, uc_1543, 
      uc_1544, uc_1545, uc_1546, uc_1547, uc_1548, uc_1549, uc_1550}), 
      .carry_final());
endmodule
