
// 	Wed Jan  4 08:21:35 2023
//	vlsi
//	192.168.44.143

module datapath__0_19 (partialProd, Acc, p_0);

output [63:0] p_0;
input [63:0] Acc;
input [63:0] partialProd;
wire n_0;
wire n_2;
wire n_1;
wire n_6;
wire n_5;
wire n_10;
wire n_9;
wire n_14;
wire n_13;
wire n_18;
wire n_17;
wire n_22;
wire n_21;
wire n_26;
wire n_25;
wire n_30;
wire n_29;
wire n_34;
wire n_33;
wire n_38;
wire n_37;
wire n_42;
wire n_41;
wire n_46;
wire n_45;
wire n_50;
wire n_49;
wire n_54;
wire n_53;
wire n_58;
wire n_57;
wire n_62;
wire n_61;
wire n_66;
wire n_65;
wire n_70;
wire n_69;
wire n_74;
wire n_73;
wire n_78;
wire n_77;
wire n_82;
wire n_81;
wire n_86;
wire n_85;
wire n_90;
wire n_89;
wire n_94;
wire n_93;
wire n_98;
wire n_97;
wire n_102;
wire n_101;
wire n_106;
wire n_105;
wire n_110;
wire n_109;
wire n_114;
wire n_113;
wire n_118;
wire n_117;
wire n_122;
wire n_121;
wire n_126;
wire n_125;
wire n_130;
wire n_129;
wire n_134;
wire n_133;
wire n_138;
wire n_137;
wire n_142;
wire n_141;
wire n_146;
wire n_145;
wire n_150;
wire n_149;
wire n_154;
wire n_153;
wire n_158;
wire n_157;
wire n_162;
wire n_161;
wire n_166;
wire n_165;
wire n_170;
wire n_169;
wire n_174;
wire n_173;
wire n_178;
wire n_177;
wire n_182;
wire n_181;
wire n_186;
wire n_185;
wire n_190;
wire n_189;
wire n_194;
wire n_193;
wire n_198;
wire n_197;
wire n_202;
wire n_201;
wire n_206;
wire n_205;
wire n_210;
wire n_209;
wire n_214;
wire n_213;
wire n_218;
wire n_217;
wire n_222;
wire n_221;
wire n_226;
wire n_225;
wire n_230;
wire n_229;
wire n_234;
wire n_233;
wire n_238;
wire n_237;
wire n_242;
wire n_241;
wire n_246;
wire n_245;
wire n_248;
wire n_244;
wire n_240;
wire n_236;
wire n_232;
wire n_228;
wire n_224;
wire n_220;
wire n_216;
wire n_212;
wire n_208;
wire n_204;
wire n_200;
wire n_196;
wire n_192;
wire n_188;
wire n_184;
wire n_180;
wire n_176;
wire n_172;
wire n_168;
wire n_164;
wire n_160;
wire n_156;
wire n_152;
wire n_148;
wire n_144;
wire n_140;
wire n_136;
wire n_132;
wire n_128;
wire n_124;
wire n_120;
wire n_116;
wire n_112;
wire n_108;
wire n_104;
wire n_100;
wire n_96;
wire n_92;
wire n_88;
wire n_84;
wire n_80;
wire n_76;
wire n_72;
wire n_68;
wire n_64;
wire n_60;
wire n_56;
wire n_52;
wire n_48;
wire n_44;
wire n_40;
wire n_36;
wire n_32;
wire n_28;
wire n_24;
wire n_20;
wire n_16;
wire n_12;
wire n_8;
wire n_4;
wire n_3;
wire n_7;
wire n_11;
wire n_15;
wire n_19;
wire n_23;
wire n_27;
wire n_31;
wire n_35;
wire n_39;
wire n_43;
wire n_47;
wire n_51;
wire n_55;
wire n_59;
wire n_63;
wire n_67;
wire n_71;
wire n_75;
wire n_79;
wire n_83;
wire n_87;
wire n_91;
wire n_95;
wire n_99;
wire n_103;
wire n_107;
wire n_111;
wire n_115;
wire n_119;
wire n_123;
wire n_127;
wire n_131;
wire n_135;
wire n_139;
wire n_143;
wire n_147;
wire n_151;
wire n_155;
wire n_159;
wire n_163;
wire n_167;
wire n_171;
wire n_175;
wire n_179;
wire n_183;
wire n_187;
wire n_191;
wire n_195;
wire n_199;
wire n_203;
wire n_207;
wire n_211;
wire n_215;
wire n_219;
wire n_223;
wire n_227;
wire n_231;
wire n_235;
wire n_239;
wire n_243;
wire n_247;


AOI21_X1 i_249 (.ZN (n_248), .A (n_2), .B1 (n_0), .B2 (n_1));
INV_X1 i_248 (.ZN (n_247), .A (n_248));
AOI21_X1 i_247 (.ZN (n_244), .A (n_6), .B1 (n_5), .B2 (n_247));
INV_X1 i_246 (.ZN (n_243), .A (n_244));
AOI21_X1 i_244 (.ZN (n_240), .A (n_10), .B1 (n_9), .B2 (n_243));
INV_X1 i_243 (.ZN (n_239), .A (n_240));
AOI21_X1 i_242 (.ZN (n_236), .A (n_14), .B1 (n_13), .B2 (n_239));
INV_X1 i_240 (.ZN (n_235), .A (n_236));
AOI21_X1 i_239 (.ZN (n_232), .A (n_18), .B1 (n_17), .B2 (n_235));
INV_X1 i_238 (.ZN (n_231), .A (n_232));
AOI21_X1 i_236 (.ZN (n_228), .A (n_22), .B1 (n_21), .B2 (n_231));
INV_X1 i_235 (.ZN (n_227), .A (n_228));
AOI21_X1 i_234 (.ZN (n_224), .A (n_26), .B1 (n_25), .B2 (n_227));
INV_X1 i_232 (.ZN (n_223), .A (n_224));
AOI21_X1 i_231 (.ZN (n_220), .A (n_30), .B1 (n_29), .B2 (n_223));
INV_X1 i_230 (.ZN (n_219), .A (n_220));
AOI21_X1 i_228 (.ZN (n_216), .A (n_34), .B1 (n_33), .B2 (n_219));
INV_X1 i_227 (.ZN (n_215), .A (n_216));
AOI21_X1 i_226 (.ZN (n_212), .A (n_38), .B1 (n_37), .B2 (n_215));
INV_X1 i_224 (.ZN (n_211), .A (n_212));
AOI21_X1 i_223 (.ZN (n_208), .A (n_42), .B1 (n_41), .B2 (n_211));
INV_X1 i_222 (.ZN (n_207), .A (n_208));
AOI21_X1 i_220 (.ZN (n_204), .A (n_46), .B1 (n_45), .B2 (n_207));
INV_X1 i_219 (.ZN (n_203), .A (n_204));
AOI21_X1 i_218 (.ZN (n_200), .A (n_50), .B1 (n_49), .B2 (n_203));
INV_X1 i_216 (.ZN (n_199), .A (n_200));
AOI21_X1 i_215 (.ZN (n_196), .A (n_54), .B1 (n_53), .B2 (n_199));
INV_X1 i_214 (.ZN (n_195), .A (n_196));
AOI21_X1 i_212 (.ZN (n_192), .A (n_58), .B1 (n_57), .B2 (n_195));
INV_X1 i_211 (.ZN (n_191), .A (n_192));
AOI21_X1 i_210 (.ZN (n_188), .A (n_62), .B1 (n_61), .B2 (n_191));
INV_X1 i_208 (.ZN (n_187), .A (n_188));
AOI21_X1 i_207 (.ZN (n_184), .A (n_66), .B1 (n_65), .B2 (n_187));
INV_X1 i_206 (.ZN (n_183), .A (n_184));
AOI21_X1 i_204 (.ZN (n_180), .A (n_70), .B1 (n_69), .B2 (n_183));
INV_X1 i_203 (.ZN (n_179), .A (n_180));
AOI21_X1 i_202 (.ZN (n_176), .A (n_74), .B1 (n_73), .B2 (n_179));
INV_X1 i_200 (.ZN (n_175), .A (n_176));
AOI21_X1 i_199 (.ZN (n_172), .A (n_78), .B1 (n_77), .B2 (n_175));
INV_X1 i_198 (.ZN (n_171), .A (n_172));
AOI21_X1 i_196 (.ZN (n_168), .A (n_82), .B1 (n_81), .B2 (n_171));
INV_X1 i_195 (.ZN (n_167), .A (n_168));
AOI21_X1 i_194 (.ZN (n_164), .A (n_86), .B1 (n_85), .B2 (n_167));
INV_X1 i_192 (.ZN (n_163), .A (n_164));
AOI21_X1 i_191 (.ZN (n_160), .A (n_90), .B1 (n_89), .B2 (n_163));
INV_X1 i_190 (.ZN (n_159), .A (n_160));
AOI21_X1 i_188 (.ZN (n_156), .A (n_94), .B1 (n_93), .B2 (n_159));
INV_X1 i_187 (.ZN (n_155), .A (n_156));
AOI21_X1 i_186 (.ZN (n_152), .A (n_98), .B1 (n_97), .B2 (n_155));
INV_X1 i_184 (.ZN (n_151), .A (n_152));
AOI21_X1 i_183 (.ZN (n_148), .A (n_102), .B1 (n_101), .B2 (n_151));
INV_X1 i_182 (.ZN (n_147), .A (n_148));
AOI21_X1 i_180 (.ZN (n_144), .A (n_106), .B1 (n_105), .B2 (n_147));
INV_X1 i_179 (.ZN (n_143), .A (n_144));
AOI21_X1 i_178 (.ZN (n_140), .A (n_110), .B1 (n_109), .B2 (n_143));
INV_X1 i_176 (.ZN (n_139), .A (n_140));
AOI21_X1 i_175 (.ZN (n_136), .A (n_114), .B1 (n_113), .B2 (n_139));
INV_X1 i_174 (.ZN (n_135), .A (n_136));
AOI21_X1 i_172 (.ZN (n_132), .A (n_118), .B1 (n_117), .B2 (n_135));
INV_X1 i_171 (.ZN (n_131), .A (n_132));
AOI21_X1 i_170 (.ZN (n_128), .A (n_122), .B1 (n_121), .B2 (n_131));
INV_X1 i_168 (.ZN (n_127), .A (n_128));
AOI21_X1 i_167 (.ZN (n_124), .A (n_126), .B1 (n_125), .B2 (n_127));
INV_X1 i_166 (.ZN (n_123), .A (n_124));
AOI21_X1 i_164 (.ZN (n_120), .A (n_130), .B1 (n_129), .B2 (n_123));
INV_X1 i_163 (.ZN (n_119), .A (n_120));
AOI21_X1 i_162 (.ZN (n_116), .A (n_134), .B1 (n_133), .B2 (n_119));
INV_X1 i_160 (.ZN (n_115), .A (n_116));
AOI21_X1 i_159 (.ZN (n_112), .A (n_138), .B1 (n_137), .B2 (n_115));
INV_X1 i_158 (.ZN (n_111), .A (n_112));
AOI21_X1 i_156 (.ZN (n_108), .A (n_142), .B1 (n_141), .B2 (n_111));
INV_X1 i_155 (.ZN (n_107), .A (n_108));
AOI21_X1 i_154 (.ZN (n_104), .A (n_146), .B1 (n_145), .B2 (n_107));
INV_X1 i_152 (.ZN (n_103), .A (n_104));
AOI21_X1 i_151 (.ZN (n_100), .A (n_150), .B1 (n_149), .B2 (n_103));
INV_X1 i_150 (.ZN (n_99), .A (n_100));
AOI21_X1 i_148 (.ZN (n_96), .A (n_154), .B1 (n_153), .B2 (n_99));
INV_X1 i_147 (.ZN (n_95), .A (n_96));
AOI21_X1 i_146 (.ZN (n_92), .A (n_158), .B1 (n_157), .B2 (n_95));
INV_X1 i_144 (.ZN (n_91), .A (n_92));
AOI21_X1 i_143 (.ZN (n_88), .A (n_162), .B1 (n_161), .B2 (n_91));
INV_X1 i_142 (.ZN (n_87), .A (n_88));
AOI21_X1 i_140 (.ZN (n_84), .A (n_166), .B1 (n_165), .B2 (n_87));
INV_X1 i_139 (.ZN (n_83), .A (n_84));
AOI21_X1 i_138 (.ZN (n_80), .A (n_170), .B1 (n_169), .B2 (n_83));
INV_X1 i_136 (.ZN (n_79), .A (n_80));
AOI21_X1 i_135 (.ZN (n_76), .A (n_174), .B1 (n_173), .B2 (n_79));
INV_X1 i_134 (.ZN (n_75), .A (n_76));
AOI21_X1 i_132 (.ZN (n_72), .A (n_178), .B1 (n_177), .B2 (n_75));
INV_X1 i_131 (.ZN (n_71), .A (n_72));
AOI21_X1 i_130 (.ZN (n_68), .A (n_182), .B1 (n_181), .B2 (n_71));
INV_X1 i_128 (.ZN (n_67), .A (n_68));
AOI21_X1 i_127 (.ZN (n_64), .A (n_186), .B1 (n_185), .B2 (n_67));
INV_X1 i_126 (.ZN (n_63), .A (n_64));
AOI21_X1 i_124 (.ZN (n_60), .A (n_190), .B1 (n_189), .B2 (n_63));
INV_X1 i_123 (.ZN (n_59), .A (n_60));
AOI21_X1 i_122 (.ZN (n_56), .A (n_194), .B1 (n_193), .B2 (n_59));
INV_X1 i_120 (.ZN (n_55), .A (n_56));
AOI21_X1 i_119 (.ZN (n_52), .A (n_198), .B1 (n_197), .B2 (n_55));
INV_X1 i_118 (.ZN (n_51), .A (n_52));
AOI21_X1 i_116 (.ZN (n_48), .A (n_202), .B1 (n_201), .B2 (n_51));
INV_X1 i_115 (.ZN (n_47), .A (n_48));
AOI21_X1 i_114 (.ZN (n_44), .A (n_206), .B1 (n_205), .B2 (n_47));
INV_X1 i_112 (.ZN (n_43), .A (n_44));
AOI21_X1 i_111 (.ZN (n_40), .A (n_210), .B1 (n_209), .B2 (n_43));
INV_X1 i_110 (.ZN (n_39), .A (n_40));
AOI21_X1 i_108 (.ZN (n_36), .A (n_214), .B1 (n_213), .B2 (n_39));
INV_X1 i_107 (.ZN (n_35), .A (n_36));
AOI21_X1 i_106 (.ZN (n_32), .A (n_218), .B1 (n_217), .B2 (n_35));
INV_X1 i_104 (.ZN (n_31), .A (n_32));
AOI21_X1 i_103 (.ZN (n_28), .A (n_222), .B1 (n_221), .B2 (n_31));
INV_X1 i_102 (.ZN (n_27), .A (n_28));
AOI21_X1 i_100 (.ZN (n_24), .A (n_226), .B1 (n_225), .B2 (n_27));
INV_X1 i_99 (.ZN (n_23), .A (n_24));
AOI21_X1 i_98 (.ZN (n_20), .A (n_230), .B1 (n_229), .B2 (n_23));
INV_X1 i_96 (.ZN (n_19), .A (n_20));
AOI21_X1 i_95 (.ZN (n_16), .A (n_234), .B1 (n_233), .B2 (n_19));
INV_X1 i_94 (.ZN (n_15), .A (n_16));
AOI21_X1 i_92 (.ZN (n_12), .A (n_238), .B1 (n_237), .B2 (n_15));
INV_X1 i_91 (.ZN (n_11), .A (n_12));
AOI21_X1 i_90 (.ZN (n_8), .A (n_242), .B1 (n_241), .B2 (n_11));
INV_X1 i_88 (.ZN (n_7), .A (n_8));
AOI21_X1 i_87 (.ZN (n_4), .A (n_246), .B1 (n_245), .B2 (n_7));
XNOR2_X1 i_86 (.ZN (n_3), .A (partialProd[63]), .B (Acc[63]));
XOR2_X1 i_84 (.Z (p_0[63]), .A (n_4), .B (n_3));
XNOR2_X1 i_83 (.ZN (p_0[62]), .A (n_245), .B (n_8));
XNOR2_X1 i_82 (.ZN (p_0[61]), .A (n_241), .B (n_12));
XNOR2_X1 i_80 (.ZN (p_0[60]), .A (n_237), .B (n_16));
XNOR2_X1 i_79 (.ZN (p_0[59]), .A (n_233), .B (n_20));
XNOR2_X1 i_78 (.ZN (p_0[58]), .A (n_229), .B (n_24));
XNOR2_X1 i_76 (.ZN (p_0[57]), .A (n_225), .B (n_28));
XNOR2_X1 i_75 (.ZN (p_0[56]), .A (n_221), .B (n_32));
XNOR2_X1 i_74 (.ZN (p_0[55]), .A (n_217), .B (n_36));
XNOR2_X1 i_72 (.ZN (p_0[54]), .A (n_213), .B (n_40));
XNOR2_X1 i_71 (.ZN (p_0[53]), .A (n_209), .B (n_44));
XNOR2_X1 i_70 (.ZN (p_0[52]), .A (n_205), .B (n_48));
XNOR2_X1 i_68 (.ZN (p_0[51]), .A (n_201), .B (n_52));
XNOR2_X1 i_67 (.ZN (p_0[50]), .A (n_197), .B (n_56));
XNOR2_X1 i_66 (.ZN (p_0[49]), .A (n_193), .B (n_60));
XNOR2_X1 i_64 (.ZN (p_0[48]), .A (n_189), .B (n_64));
XNOR2_X1 i_63 (.ZN (p_0[47]), .A (n_185), .B (n_68));
XNOR2_X1 i_62 (.ZN (p_0[46]), .A (n_181), .B (n_72));
XNOR2_X1 i_60 (.ZN (p_0[45]), .A (n_177), .B (n_76));
XNOR2_X1 i_59 (.ZN (p_0[44]), .A (n_173), .B (n_80));
XNOR2_X1 i_58 (.ZN (p_0[43]), .A (n_169), .B (n_84));
XNOR2_X1 i_56 (.ZN (p_0[42]), .A (n_165), .B (n_88));
XNOR2_X1 i_55 (.ZN (p_0[41]), .A (n_161), .B (n_92));
XNOR2_X1 i_54 (.ZN (p_0[40]), .A (n_157), .B (n_96));
XNOR2_X1 i_52 (.ZN (p_0[39]), .A (n_153), .B (n_100));
XNOR2_X1 i_51 (.ZN (p_0[38]), .A (n_149), .B (n_104));
XNOR2_X1 i_50 (.ZN (p_0[37]), .A (n_145), .B (n_108));
XNOR2_X1 i_48 (.ZN (p_0[36]), .A (n_141), .B (n_112));
XNOR2_X1 i_47 (.ZN (p_0[35]), .A (n_137), .B (n_116));
XNOR2_X1 i_46 (.ZN (p_0[34]), .A (n_133), .B (n_120));
XNOR2_X1 i_44 (.ZN (p_0[33]), .A (n_129), .B (n_124));
XNOR2_X1 i_43 (.ZN (p_0[32]), .A (n_125), .B (n_128));
XNOR2_X1 i_42 (.ZN (p_0[31]), .A (n_121), .B (n_132));
XNOR2_X1 i_40 (.ZN (p_0[30]), .A (n_117), .B (n_136));
XNOR2_X1 i_39 (.ZN (p_0[29]), .A (n_113), .B (n_140));
XNOR2_X1 i_38 (.ZN (p_0[28]), .A (n_109), .B (n_144));
XNOR2_X1 i_36 (.ZN (p_0[27]), .A (n_105), .B (n_148));
XNOR2_X1 i_35 (.ZN (p_0[26]), .A (n_101), .B (n_152));
XNOR2_X1 i_34 (.ZN (p_0[25]), .A (n_97), .B (n_156));
XNOR2_X1 i_32 (.ZN (p_0[24]), .A (n_93), .B (n_160));
XNOR2_X1 i_31 (.ZN (p_0[23]), .A (n_89), .B (n_164));
XNOR2_X1 i_30 (.ZN (p_0[22]), .A (n_85), .B (n_168));
XNOR2_X1 i_28 (.ZN (p_0[21]), .A (n_81), .B (n_172));
XNOR2_X1 i_27 (.ZN (p_0[20]), .A (n_77), .B (n_176));
XNOR2_X1 i_26 (.ZN (p_0[19]), .A (n_73), .B (n_180));
XNOR2_X1 i_24 (.ZN (p_0[18]), .A (n_69), .B (n_184));
XNOR2_X1 i_23 (.ZN (p_0[17]), .A (n_65), .B (n_188));
XNOR2_X1 i_22 (.ZN (p_0[16]), .A (n_61), .B (n_192));
XNOR2_X1 i_20 (.ZN (p_0[15]), .A (n_57), .B (n_196));
XNOR2_X1 i_19 (.ZN (p_0[14]), .A (n_53), .B (n_200));
XNOR2_X1 i_18 (.ZN (p_0[13]), .A (n_49), .B (n_204));
XNOR2_X1 i_16 (.ZN (p_0[12]), .A (n_45), .B (n_208));
XNOR2_X1 i_15 (.ZN (p_0[11]), .A (n_41), .B (n_212));
XNOR2_X1 i_14 (.ZN (p_0[10]), .A (n_37), .B (n_216));
XNOR2_X1 i_12 (.ZN (p_0[9]), .A (n_33), .B (n_220));
XNOR2_X1 i_11 (.ZN (p_0[8]), .A (n_29), .B (n_224));
XNOR2_X1 i_10 (.ZN (p_0[7]), .A (n_25), .B (n_228));
XNOR2_X1 i_8 (.ZN (p_0[6]), .A (n_21), .B (n_232));
XNOR2_X1 i_7 (.ZN (p_0[5]), .A (n_17), .B (n_236));
XNOR2_X1 i_6 (.ZN (p_0[4]), .A (n_13), .B (n_240));
XNOR2_X1 i_4 (.ZN (p_0[3]), .A (n_9), .B (n_244));
XNOR2_X1 i_3 (.ZN (p_0[2]), .A (n_5), .B (n_248));
XOR2_X1 i_2 (.Z (p_0[1]), .A (n_0), .B (n_1));
HA_X1 i_245 (.CO (n_246), .S (n_245), .A (partialProd[62]), .B (Acc[62]));
HA_X1 i_241 (.CO (n_242), .S (n_241), .A (partialProd[61]), .B (Acc[61]));
HA_X1 i_237 (.CO (n_238), .S (n_237), .A (partialProd[60]), .B (Acc[60]));
HA_X1 i_233 (.CO (n_234), .S (n_233), .A (partialProd[59]), .B (Acc[59]));
HA_X1 i_229 (.CO (n_230), .S (n_229), .A (partialProd[58]), .B (Acc[58]));
HA_X1 i_225 (.CO (n_226), .S (n_225), .A (partialProd[57]), .B (Acc[57]));
HA_X1 i_221 (.CO (n_222), .S (n_221), .A (partialProd[56]), .B (Acc[56]));
HA_X1 i_217 (.CO (n_218), .S (n_217), .A (partialProd[55]), .B (Acc[55]));
HA_X1 i_213 (.CO (n_214), .S (n_213), .A (partialProd[54]), .B (Acc[54]));
HA_X1 i_209 (.CO (n_210), .S (n_209), .A (partialProd[53]), .B (Acc[53]));
HA_X1 i_205 (.CO (n_206), .S (n_205), .A (partialProd[52]), .B (Acc[52]));
HA_X1 i_201 (.CO (n_202), .S (n_201), .A (partialProd[51]), .B (Acc[51]));
HA_X1 i_197 (.CO (n_198), .S (n_197), .A (partialProd[50]), .B (Acc[50]));
HA_X1 i_193 (.CO (n_194), .S (n_193), .A (partialProd[49]), .B (Acc[49]));
HA_X1 i_189 (.CO (n_190), .S (n_189), .A (partialProd[48]), .B (Acc[48]));
HA_X1 i_185 (.CO (n_186), .S (n_185), .A (partialProd[47]), .B (Acc[47]));
HA_X1 i_181 (.CO (n_182), .S (n_181), .A (partialProd[46]), .B (Acc[46]));
HA_X1 i_177 (.CO (n_178), .S (n_177), .A (partialProd[45]), .B (Acc[45]));
HA_X1 i_173 (.CO (n_174), .S (n_173), .A (partialProd[44]), .B (Acc[44]));
HA_X1 i_169 (.CO (n_170), .S (n_169), .A (partialProd[43]), .B (Acc[43]));
HA_X1 i_165 (.CO (n_166), .S (n_165), .A (partialProd[42]), .B (Acc[42]));
HA_X1 i_161 (.CO (n_162), .S (n_161), .A (partialProd[41]), .B (Acc[41]));
HA_X1 i_157 (.CO (n_158), .S (n_157), .A (partialProd[40]), .B (Acc[40]));
HA_X1 i_153 (.CO (n_154), .S (n_153), .A (partialProd[39]), .B (Acc[39]));
HA_X1 i_149 (.CO (n_150), .S (n_149), .A (partialProd[38]), .B (Acc[38]));
HA_X1 i_145 (.CO (n_146), .S (n_145), .A (partialProd[37]), .B (Acc[37]));
HA_X1 i_141 (.CO (n_142), .S (n_141), .A (partialProd[36]), .B (Acc[36]));
HA_X1 i_137 (.CO (n_138), .S (n_137), .A (partialProd[35]), .B (Acc[35]));
HA_X1 i_133 (.CO (n_134), .S (n_133), .A (partialProd[34]), .B (Acc[34]));
HA_X1 i_129 (.CO (n_130), .S (n_129), .A (partialProd[33]), .B (Acc[33]));
HA_X1 i_125 (.CO (n_126), .S (n_125), .A (partialProd[32]), .B (Acc[32]));
HA_X1 i_121 (.CO (n_122), .S (n_121), .A (partialProd[31]), .B (Acc[31]));
HA_X1 i_117 (.CO (n_118), .S (n_117), .A (partialProd[30]), .B (Acc[30]));
HA_X1 i_113 (.CO (n_114), .S (n_113), .A (partialProd[29]), .B (Acc[29]));
HA_X1 i_109 (.CO (n_110), .S (n_109), .A (partialProd[28]), .B (Acc[28]));
HA_X1 i_105 (.CO (n_106), .S (n_105), .A (partialProd[27]), .B (Acc[27]));
HA_X1 i_101 (.CO (n_102), .S (n_101), .A (partialProd[26]), .B (Acc[26]));
HA_X1 i_97 (.CO (n_98), .S (n_97), .A (partialProd[25]), .B (Acc[25]));
HA_X1 i_93 (.CO (n_94), .S (n_93), .A (partialProd[24]), .B (Acc[24]));
HA_X1 i_89 (.CO (n_90), .S (n_89), .A (partialProd[23]), .B (Acc[23]));
HA_X1 i_85 (.CO (n_86), .S (n_85), .A (partialProd[22]), .B (Acc[22]));
HA_X1 i_81 (.CO (n_82), .S (n_81), .A (partialProd[21]), .B (Acc[21]));
HA_X1 i_77 (.CO (n_78), .S (n_77), .A (partialProd[20]), .B (Acc[20]));
HA_X1 i_73 (.CO (n_74), .S (n_73), .A (partialProd[19]), .B (Acc[19]));
HA_X1 i_69 (.CO (n_70), .S (n_69), .A (partialProd[18]), .B (Acc[18]));
HA_X1 i_65 (.CO (n_66), .S (n_65), .A (partialProd[17]), .B (Acc[17]));
HA_X1 i_61 (.CO (n_62), .S (n_61), .A (partialProd[16]), .B (Acc[16]));
HA_X1 i_57 (.CO (n_58), .S (n_57), .A (partialProd[15]), .B (Acc[15]));
HA_X1 i_53 (.CO (n_54), .S (n_53), .A (partialProd[14]), .B (Acc[14]));
HA_X1 i_49 (.CO (n_50), .S (n_49), .A (partialProd[13]), .B (Acc[13]));
HA_X1 i_45 (.CO (n_46), .S (n_45), .A (partialProd[12]), .B (Acc[12]));
HA_X1 i_41 (.CO (n_42), .S (n_41), .A (partialProd[11]), .B (Acc[11]));
HA_X1 i_37 (.CO (n_38), .S (n_37), .A (partialProd[10]), .B (Acc[10]));
HA_X1 i_33 (.CO (n_34), .S (n_33), .A (partialProd[9]), .B (Acc[9]));
HA_X1 i_29 (.CO (n_30), .S (n_29), .A (partialProd[8]), .B (Acc[8]));
HA_X1 i_25 (.CO (n_26), .S (n_25), .A (partialProd[7]), .B (Acc[7]));
HA_X1 i_21 (.CO (n_22), .S (n_21), .A (partialProd[6]), .B (Acc[6]));
HA_X1 i_17 (.CO (n_18), .S (n_17), .A (partialProd[5]), .B (Acc[5]));
HA_X1 i_13 (.CO (n_14), .S (n_13), .A (partialProd[4]), .B (Acc[4]));
HA_X1 i_9 (.CO (n_10), .S (n_9), .A (partialProd[3]), .B (Acc[3]));
HA_X1 i_5 (.CO (n_6), .S (n_5), .A (partialProd[2]), .B (Acc[2]));
HA_X1 i_1 (.CO (n_2), .S (n_1), .A (partialProd[1]), .B (Acc[1]));
HA_X1 i_0 (.CO (n_0), .S (p_0[0]), .A (partialProd[0]), .B (Acc[0]));

endmodule //datapath__0_19

module datapath (p_0, A_reg);

output [31:0] p_0;
input [31:0] A_reg;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (A_reg[25]));
INV_X1 i_63 (.ZN (n_32), .A (A_reg[21]));
INV_X1 i_62 (.ZN (n_31), .A (A_reg[14]));
INV_X1 i_61 (.ZN (n_30), .A (A_reg[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (A_reg[2]), .A2 (A_reg[1]), .A3 (A_reg[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (A_reg[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (A_reg[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (A_reg[5]), .A3 (A_reg[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (A_reg[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (A_reg[8]), .A3 (A_reg[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (A_reg[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (A_reg[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (A_reg[12]), .A3 (A_reg[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (A_reg[15]), .A3 (A_reg[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (A_reg[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (A_reg[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (A_reg[18]), .A3 (A_reg[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (A_reg[18]), .A3 (A_reg[19]), .A4 (A_reg[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (A_reg[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (A_reg[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (A_reg[23]), .A3 (A_reg[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (A_reg[26]), .A3 (A_reg[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (A_reg[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (A_reg[28]), .A3 (A_reg[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (A_reg[28]), .A3 (A_reg[29]), .A4 (A_reg[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (A_reg[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (A_reg[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (A_reg[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (A_reg[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (A_reg[27]), .B1 (n_9), .B2 (A_reg[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (A_reg[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (A_reg[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (A_reg[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (A_reg[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (A_reg[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (A_reg[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (A_reg[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (A_reg[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (A_reg[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (A_reg[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (A_reg[16]), .B1 (n_19), .B2 (A_reg[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (A_reg[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (A_reg[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (A_reg[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (A_reg[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (A_reg[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (A_reg[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (A_reg[9]), .B1 (n_25), .B2 (A_reg[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (A_reg[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (A_reg[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (A_reg[6]), .B1 (n_27), .B2 (A_reg[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (A_reg[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (A_reg[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (A_reg[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (A_reg[2]), .B1 (A_reg[1]), .B2 (A_reg[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (A_reg[1]), .B (A_reg[0]));

endmodule //datapath

module registerNbits__parameterized0 (clk_CTSPP_1, clk, reset, en, inp, out);

output [63:0] out;
input clk;
input en;
input [63:0] inp;
input reset;
input clk_CTSPP_1;
wire n_0_0;
wire n_1;
wire CTS_n10;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire hfn_ipo_n5;
wire CTS_n11;


AND2_X1 i_0_65 (.ZN (n_65), .A1 (hfn_ipo_n5), .A2 (inp[63]));
AND2_X1 i_0_64 (.ZN (n_64), .A1 (hfn_ipo_n5), .A2 (inp[62]));
AND2_X1 i_0_63 (.ZN (n_63), .A1 (hfn_ipo_n5), .A2 (inp[61]));
AND2_X1 i_0_62 (.ZN (n_62), .A1 (hfn_ipo_n5), .A2 (inp[60]));
AND2_X1 i_0_61 (.ZN (n_61), .A1 (hfn_ipo_n5), .A2 (inp[59]));
AND2_X1 i_0_60 (.ZN (n_60), .A1 (hfn_ipo_n5), .A2 (inp[58]));
AND2_X1 i_0_59 (.ZN (n_59), .A1 (hfn_ipo_n5), .A2 (inp[57]));
AND2_X1 i_0_58 (.ZN (n_58), .A1 (hfn_ipo_n5), .A2 (inp[56]));
AND2_X1 i_0_57 (.ZN (n_57), .A1 (hfn_ipo_n5), .A2 (inp[55]));
AND2_X1 i_0_56 (.ZN (n_56), .A1 (hfn_ipo_n5), .A2 (inp[54]));
AND2_X1 i_0_55 (.ZN (n_55), .A1 (hfn_ipo_n5), .A2 (inp[53]));
AND2_X1 i_0_54 (.ZN (n_54), .A1 (hfn_ipo_n5), .A2 (inp[52]));
AND2_X1 i_0_53 (.ZN (n_53), .A1 (hfn_ipo_n5), .A2 (inp[51]));
AND2_X1 i_0_52 (.ZN (n_52), .A1 (hfn_ipo_n5), .A2 (inp[50]));
AND2_X1 i_0_51 (.ZN (n_51), .A1 (hfn_ipo_n5), .A2 (inp[49]));
AND2_X1 i_0_50 (.ZN (n_50), .A1 (hfn_ipo_n5), .A2 (inp[48]));
AND2_X1 i_0_49 (.ZN (n_49), .A1 (hfn_ipo_n5), .A2 (inp[47]));
AND2_X1 i_0_48 (.ZN (n_48), .A1 (hfn_ipo_n5), .A2 (inp[46]));
AND2_X1 i_0_47 (.ZN (n_47), .A1 (hfn_ipo_n5), .A2 (inp[45]));
AND2_X1 i_0_46 (.ZN (n_46), .A1 (hfn_ipo_n5), .A2 (inp[44]));
AND2_X1 i_0_45 (.ZN (n_45), .A1 (hfn_ipo_n5), .A2 (inp[43]));
AND2_X1 i_0_44 (.ZN (n_44), .A1 (hfn_ipo_n5), .A2 (inp[42]));
AND2_X1 i_0_43 (.ZN (n_43), .A1 (hfn_ipo_n5), .A2 (inp[41]));
AND2_X1 i_0_42 (.ZN (n_42), .A1 (hfn_ipo_n5), .A2 (inp[40]));
AND2_X1 i_0_41 (.ZN (n_41), .A1 (n_0_0), .A2 (inp[39]));
AND2_X1 i_0_40 (.ZN (n_40), .A1 (n_0_0), .A2 (inp[38]));
AND2_X1 i_0_39 (.ZN (n_39), .A1 (n_0_0), .A2 (inp[37]));
AND2_X1 i_0_38 (.ZN (n_38), .A1 (n_0_0), .A2 (inp[36]));
AND2_X1 i_0_37 (.ZN (n_37), .A1 (n_0_0), .A2 (inp[35]));
AND2_X1 i_0_36 (.ZN (n_36), .A1 (n_0_0), .A2 (inp[34]));
AND2_X1 i_0_35 (.ZN (n_35), .A1 (n_0_0), .A2 (inp[33]));
AND2_X1 i_0_34 (.ZN (n_34), .A1 (n_0_0), .A2 (inp[32]));
AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (hfn_ipo_n5), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (hfn_ipo_n5), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (hfn_ipo_n5), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (hfn_ipo_n5), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (hfn_ipo_n5), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (hfn_ipo_n5), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (hfn_ipo_n5), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (hfn_ipo_n5), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (hfn_ipo_n5), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (hfn_ipo_n5), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (hfn_ipo_n5), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (hfn_ipo_n5), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (hfn_ipo_n5), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (hfn_ipo_n5), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (hfn_ipo_n5), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n10), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n10), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n10), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n10), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n10), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n10), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n10), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n10), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n10), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n10), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n10), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n10), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n10), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n10), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n10), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n10), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n10), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n10), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n10), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n10), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n10), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n10), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n10), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n10), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n10), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n10), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n10), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n10), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n10), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n10), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n10), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n10), .D (n_33));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (CTS_n10), .D (n_34));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (CTS_n10), .D (n_35));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (CTS_n10), .D (n_36));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (CTS_n10), .D (n_37));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (CTS_n10), .D (n_38));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (CTS_n10), .D (n_39));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (CTS_n10), .D (n_40));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (CTS_n10), .D (n_41));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (CTS_n10), .D (n_42));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (CTS_n10), .D (n_43));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (CTS_n10), .D (n_44));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (CTS_n10), .D (n_45));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (CTS_n10), .D (n_46));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (CTS_n10), .D (n_47));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (CTS_n10), .D (n_48));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (CTS_n10), .D (n_49));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (CTS_n10), .D (n_50));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (CTS_n10), .D (n_51));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (CTS_n10), .D (n_52));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (CTS_n10), .D (n_53));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (CTS_n10), .D (n_54));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (CTS_n10), .D (n_55));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (CTS_n10), .D (n_56));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (CTS_n10), .D (n_57));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (CTS_n10), .D (n_58));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (CTS_n10), .D (n_59));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (CTS_n10), .D (n_60));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (CTS_n10), .D (n_61));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (CTS_n10), .D (n_62));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (CTS_n10), .D (n_63));
DFF_X1 \out_reg[62]  (.Q (out[62]), .CK (CTS_n10), .D (n_64));
DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (CTS_n10), .D (n_65));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n11), .CK (clk_CTSPP_1), .E (n_1), .SE (VSS));
BUF_X4 hfn_ipo_c5 (.Z (hfn_ipo_n5), .A (n_0_0));
CLKBUF_X3 CTS_L3_c11 (.Z (CTS_n10), .A (CTS_n11));

endmodule //registerNbits__parameterized0

module registerNbits (clk_CTSPP_1, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTSPP_1;
wire CLOCK_slh__n23;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CLOCK_slh__n25;
wire CLOCK_slh__n27;
wire CLOCK_slh__n29;
wire CLOCK_slh__n31;
wire CLOCK_slh__n33;
wire CLOCK_slh__n35;
wire CLOCK_slh__n37;
wire CLOCK_slh__n39;
wire CLOCK_slh__n41;
wire CLOCK_slh__n43;
wire CLOCK_slh__n45;
wire CLOCK_slh__n47;
wire CLOCK_slh__n49;
wire CLOCK_slh__n51;
wire CLOCK_slh__n53;
wire CLOCK_slh__n55;
wire CLOCK_slh__n57;
wire CLOCK_slh__n59;
wire CLOCK_slh__n61;
wire CLOCK_slh__n63;
wire CLOCK_slh__n65;
wire CLOCK_slh__n67;
wire CLOCK_slh__n69;
wire CLOCK_slh__n71;
wire CLOCK_slh__n73;
wire CLOCK_slh__n75;
wire CLOCK_slh__n77;
wire CLOCK_slh__n79;
wire CLOCK_slh__n81;
wire CLOCK_slh__n83;
wire CLOCK_slh__n85;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n25), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n23), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n59), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n35), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n37), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n33), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n41), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n71), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n75), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n69), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n57), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n85), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n51), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n63), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n83), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n77), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n73), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n65), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n39), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n61), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n67), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n49), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n27), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n55), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n81), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n47), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n79), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n53), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n31), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n29), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n45), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n43), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTSPP_1), .E (n_1), .SE (VSS));
CLKBUF_X1 CLOCK_slh__c7 (.Z (n_32), .A (CLOCK_slh__n23));
CLKBUF_X1 CLOCK_slh__c9 (.Z (n_33), .A (CLOCK_slh__n25));
CLKBUF_X1 CLOCK_slh__c11 (.Z (n_11), .A (CLOCK_slh__n27));
CLKBUF_X1 CLOCK_slh__c13 (.Z (n_4), .A (CLOCK_slh__n29));
CLKBUF_X1 CLOCK_slh__c15 (.Z (n_5), .A (CLOCK_slh__n31));
CLKBUF_X1 CLOCK_slh__c17 (.Z (n_28), .A (CLOCK_slh__n33));
CLKBUF_X1 CLOCK_slh__c19 (.Z (n_30), .A (CLOCK_slh__n35));
CLKBUF_X1 CLOCK_slh__c21 (.Z (n_29), .A (CLOCK_slh__n37));
CLKBUF_X1 CLOCK_slh__c23 (.Z (n_15), .A (CLOCK_slh__n39));
CLKBUF_X1 CLOCK_slh__c25 (.Z (n_27), .A (CLOCK_slh__n41));
CLKBUF_X1 CLOCK_slh__c27 (.Z (n_2), .A (CLOCK_slh__n43));
CLKBUF_X1 CLOCK_slh__c29 (.Z (n_3), .A (CLOCK_slh__n45));
CLKBUF_X1 CLOCK_slh__c31 (.Z (n_8), .A (CLOCK_slh__n47));
CLKBUF_X1 CLOCK_slh__c33 (.Z (n_12), .A (CLOCK_slh__n49));
CLKBUF_X1 CLOCK_slh__c35 (.Z (n_21), .A (CLOCK_slh__n51));
CLKBUF_X1 CLOCK_slh__c37 (.Z (n_6), .A (CLOCK_slh__n53));
CLKBUF_X1 CLOCK_slh__c39 (.Z (n_10), .A (CLOCK_slh__n55));
CLKBUF_X1 CLOCK_slh__c41 (.Z (n_23), .A (CLOCK_slh__n57));
CLKBUF_X1 CLOCK_slh__c43 (.Z (n_31), .A (CLOCK_slh__n59));
CLKBUF_X1 CLOCK_slh__c45 (.Z (n_14), .A (CLOCK_slh__n61));
CLKBUF_X1 CLOCK_slh__c47 (.Z (n_20), .A (CLOCK_slh__n63));
CLKBUF_X1 CLOCK_slh__c49 (.Z (n_16), .A (CLOCK_slh__n65));
CLKBUF_X1 CLOCK_slh__c51 (.Z (n_13), .A (CLOCK_slh__n67));
CLKBUF_X1 CLOCK_slh__c53 (.Z (n_24), .A (CLOCK_slh__n69));
CLKBUF_X1 CLOCK_slh__c55 (.Z (n_26), .A (CLOCK_slh__n71));
CLKBUF_X1 CLOCK_slh__c57 (.Z (n_17), .A (CLOCK_slh__n73));
CLKBUF_X1 CLOCK_slh__c59 (.Z (n_25), .A (CLOCK_slh__n75));
CLKBUF_X1 CLOCK_slh__c61 (.Z (n_18), .A (CLOCK_slh__n77));
CLKBUF_X1 CLOCK_slh__c63 (.Z (n_7), .A (CLOCK_slh__n79));
CLKBUF_X1 CLOCK_slh__c65 (.Z (n_9), .A (CLOCK_slh__n81));
CLKBUF_X1 CLOCK_slh__c67 (.Z (n_19), .A (CLOCK_slh__n83));
CLKBUF_X1 CLOCK_slh__c69 (.Z (n_22), .A (CLOCK_slh__n85));

endmodule //registerNbits

module registerNbits__0_23 (clk_CTSPP_1, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTSPP_1;
wire CLOCK_slh__n23;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CLOCK_slh__n25;
wire CLOCK_slh__n27;
wire CLOCK_slh__n29;
wire CLOCK_slh__n31;
wire CLOCK_slh__n33;
wire CLOCK_slh__n35;
wire CLOCK_slh__n37;
wire CLOCK_slh__n39;
wire CLOCK_slh__n41;
wire CLOCK_slh__n43;
wire CLOCK_slh__n45;
wire CLOCK_slh__n47;
wire CLOCK_slh__n49;
wire CLOCK_slh__n51;
wire CLOCK_slh__n53;
wire CLOCK_slh__n55;
wire CLOCK_slh__n57;
wire CLOCK_slh__n59;
wire CLOCK_slh__n61;
wire CLOCK_slh__n63;
wire CLOCK_slh__n65;
wire CLOCK_slh__n67;
wire CLOCK_slh__n69;
wire CLOCK_slh__n71;
wire CLOCK_slh__n73;
wire CLOCK_slh__n75;
wire CLOCK_slh__n77;
wire CLOCK_slh__n79;
wire CLOCK_slh__n81;
wire CLOCK_slh__n83;
wire CLOCK_slh__n85;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n45), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n85), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n51), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n41), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n37), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n77), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n23), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n81), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n35), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n57), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n33), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n31), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n53), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n73), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n61), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n79), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n49), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n59), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n71), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n29), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n27), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n75), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n25), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n63), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n43), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n69), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n55), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n67), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n47), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n83), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n39), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n65), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTSPP_1), .E (n_1), .SE (VSS));
CLKBUF_X1 CLOCK_slh__c7 (.Z (n_27), .A (CLOCK_slh__n23));
CLKBUF_X1 CLOCK_slh__c9 (.Z (n_11), .A (CLOCK_slh__n25));
CLKBUF_X1 CLOCK_slh__c11 (.Z (n_13), .A (CLOCK_slh__n27));
CLKBUF_X1 CLOCK_slh__c13 (.Z (n_14), .A (CLOCK_slh__n29));
CLKBUF_X1 CLOCK_slh__c15 (.Z (n_22), .A (CLOCK_slh__n31));
CLKBUF_X1 CLOCK_slh__c17 (.Z (n_23), .A (CLOCK_slh__n33));
CLKBUF_X1 CLOCK_slh__c19 (.Z (n_25), .A (CLOCK_slh__n35));
CLKBUF_X1 CLOCK_slh__c21 (.Z (n_29), .A (CLOCK_slh__n37));
CLKBUF_X1 CLOCK_slh__c23 (.Z (n_3), .A (CLOCK_slh__n39));
CLKBUF_X1 CLOCK_slh__c25 (.Z (n_30), .A (CLOCK_slh__n41));
CLKBUF_X1 CLOCK_slh__c27 (.Z (n_9), .A (CLOCK_slh__n43));
CLKBUF_X1 CLOCK_slh__c29 (.Z (n_33), .A (CLOCK_slh__n45));
CLKBUF_X1 CLOCK_slh__c31 (.Z (n_5), .A (CLOCK_slh__n47));
CLKBUF_X1 CLOCK_slh__c33 (.Z (n_17), .A (CLOCK_slh__n49));
CLKBUF_X1 CLOCK_slh__c35 (.Z (n_31), .A (CLOCK_slh__n51));
CLKBUF_X1 CLOCK_slh__c37 (.Z (n_21), .A (CLOCK_slh__n53));
CLKBUF_X1 CLOCK_slh__c39 (.Z (n_7), .A (CLOCK_slh__n55));
CLKBUF_X1 CLOCK_slh__c41 (.Z (n_24), .A (CLOCK_slh__n57));
CLKBUF_X1 CLOCK_slh__c43 (.Z (n_16), .A (CLOCK_slh__n59));
CLKBUF_X1 CLOCK_slh__c45 (.Z (n_19), .A (CLOCK_slh__n61));
CLKBUF_X1 CLOCK_slh__c47 (.Z (n_10), .A (CLOCK_slh__n63));
CLKBUF_X1 CLOCK_slh__c49 (.Z (n_2), .A (CLOCK_slh__n65));
CLKBUF_X1 CLOCK_slh__c51 (.Z (n_6), .A (CLOCK_slh__n67));
CLKBUF_X1 CLOCK_slh__c53 (.Z (n_8), .A (CLOCK_slh__n69));
CLKBUF_X1 CLOCK_slh__c55 (.Z (n_15), .A (CLOCK_slh__n71));
CLKBUF_X1 CLOCK_slh__c57 (.Z (n_20), .A (CLOCK_slh__n73));
CLKBUF_X1 CLOCK_slh__c59 (.Z (n_12), .A (CLOCK_slh__n75));
CLKBUF_X1 CLOCK_slh__c61 (.Z (n_28), .A (CLOCK_slh__n77));
CLKBUF_X1 CLOCK_slh__c63 (.Z (n_18), .A (CLOCK_slh__n79));
CLKBUF_X1 CLOCK_slh__c65 (.Z (n_26), .A (CLOCK_slh__n81));
CLKBUF_X1 CLOCK_slh__c67 (.Z (n_4), .A (CLOCK_slh__n83));
CLKBUF_X1 CLOCK_slh__c69 (.Z (n_32), .A (CLOCK_slh__n85));

endmodule //registerNbits__0_23

module RadixBooth (inputA, inputB, result, clk, reset, en, start);

output [63:0] result;
input clk;
input en;
input [31:0] inputA;
input [31:0] inputB;
input reset;
input start;
wire CLOCK_slh_n317;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire CTS_n214;
wire \out_reg[63] ;
wire \out_reg[62] ;
wire \out_reg[61] ;
wire \out_reg[60] ;
wire \out_reg[59] ;
wire \out_reg[58] ;
wire \out_reg[57] ;
wire \out_reg[56] ;
wire \out_reg[55] ;
wire \out_reg[54] ;
wire \out_reg[53] ;
wire \out_reg[52] ;
wire \out_reg[51] ;
wire \out_reg[50] ;
wire \out_reg[49] ;
wire \out_reg[48] ;
wire \out_reg[47] ;
wire \out_reg[46] ;
wire \out_reg[45] ;
wire \out_reg[44] ;
wire \out_reg[43] ;
wire \out_reg[42] ;
wire \out_reg[41] ;
wire \out_reg[40] ;
wire \out_reg[39] ;
wire \out_reg[38] ;
wire \out_reg[37] ;
wire \out_reg[36] ;
wire \out_reg[35] ;
wire \out_reg[34] ;
wire \out_reg[33] ;
wire \out_reg[32] ;
wire \out_reg[31] ;
wire \out_reg[30] ;
wire \out_reg[29] ;
wire \out_reg[28] ;
wire \out_reg[27] ;
wire \out_reg[26] ;
wire \out_reg[25] ;
wire \out_reg[24] ;
wire \out_reg[23] ;
wire \out_reg[22] ;
wire \out_reg[21] ;
wire \out_reg[20] ;
wire \out_reg[19] ;
wire \out_reg[18] ;
wire \out_reg[17] ;
wire \out_reg[16] ;
wire \out_reg[15] ;
wire \out_reg[14] ;
wire \out_reg[13] ;
wire \out_reg[12] ;
wire \out_reg[11] ;
wire \out_reg[10] ;
wire \out_reg[9] ;
wire \out_reg[8] ;
wire \out_reg[7] ;
wire \out_reg[6] ;
wire \out_reg[5] ;
wire \out_reg[4] ;
wire \out_reg[3] ;
wire \out_reg[2] ;
wire \out_reg[1] ;
wire \out_reg[0] ;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_1;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_78;
wire n_0_79;
wire n_0_80;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_0_3;
wire n_0_0_0;
wire n_0_0_4;
wire n_0_0_1;
wire n_0_0_5;
wire n_0_0_2;
wire n_0_0_6;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_0_39;
wire n_0_0_40;
wire n_0_0_41;
wire n_0_0_42;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire n_0_0_47;
wire n_0_0_48;
wire n_0_0_49;
wire n_0_0_50;
wire n_0_0_51;
wire n_0_0_52;
wire n_0_0_53;
wire n_0_0_54;
wire n_0_0_55;
wire n_0_0_56;
wire n_0_0_57;
wire n_0_0_58;
wire n_0_0_59;
wire \partialProd[63] ;
wire \partialProd[62] ;
wire \partialProd[61] ;
wire \partialProd[60] ;
wire \partialProd[59] ;
wire \partialProd[58] ;
wire \partialProd[57] ;
wire \partialProd[56] ;
wire \partialProd[55] ;
wire \partialProd[54] ;
wire \partialProd[53] ;
wire \partialProd[52] ;
wire \partialProd[51] ;
wire \partialProd[50] ;
wire \partialProd[49] ;
wire \partialProd[48] ;
wire \partialProd[47] ;
wire \partialProd[46] ;
wire \partialProd[45] ;
wire \partialProd[44] ;
wire \partialProd[43] ;
wire \partialProd[42] ;
wire \partialProd[41] ;
wire \partialProd[40] ;
wire \partialProd[39] ;
wire \partialProd[38] ;
wire \partialProd[37] ;
wire \partialProd[36] ;
wire \partialProd[35] ;
wire \partialProd[34] ;
wire \partialProd[33] ;
wire \partialProd[32] ;
wire \partialProd[31] ;
wire \partialProd[30] ;
wire \partialProd[29] ;
wire \partialProd[28] ;
wire \partialProd[27] ;
wire \partialProd[26] ;
wire \partialProd[25] ;
wire \partialProd[24] ;
wire \partialProd[23] ;
wire \partialProd[22] ;
wire \partialProd[21] ;
wire \partialProd[20] ;
wire \partialProd[19] ;
wire \partialProd[18] ;
wire \partialProd[17] ;
wire \partialProd[16] ;
wire \partialProd[15] ;
wire \partialProd[14] ;
wire \partialProd[13] ;
wire \partialProd[12] ;
wire \partialProd[11] ;
wire \partialProd[10] ;
wire \partialProd[9] ;
wire \partialProd[8] ;
wire \partialProd[7] ;
wire \partialProd[6] ;
wire \partialProd[5] ;
wire \partialProd[4] ;
wire \partialProd[3] ;
wire \partialProd[2] ;
wire \partialProd[1] ;
wire \partialProd[0] ;
wire n_0_0_60;
wire n_0_0_61;
wire n_0_0_62;
wire n_0_0_63;
wire n_0_0_64;
wire n_0_0_65;
wire n_0_0_66;
wire n_0_0_67;
wire n_0_0_68;
wire n_0_0_69;
wire n_0_0_70;
wire n_0_0_71;
wire n_0_0_72;
wire n_0_0_73;
wire n_0_0_74;
wire n_0_0_75;
wire n_0_0_76;
wire n_0_0_77;
wire n_0_0_78;
wire n_0_0_79;
wire n_0_0_80;
wire n_0_0_81;
wire n_0_0_82;
wire n_0_0_83;
wire n_0_0_84;
wire n_0_0_85;
wire n_0_0_86;
wire n_0_0_87;
wire n_0_0_88;
wire n_0_0_89;
wire n_0_0_90;
wire n_0_0_91;
wire n_0_0_92;
wire n_0_0_93;
wire n_0_0_94;
wire n_0_0_95;
wire n_0_0_96;
wire n_0_0_97;
wire n_0_0_98;
wire n_0_0_99;
wire n_0_0_100;
wire n_0_0_101;
wire n_0_0_102;
wire n_0_0_103;
wire n_0_0_104;
wire n_0_0_105;
wire n_0_0_106;
wire n_0_0_107;
wire n_0_0_108;
wire n_0_0_109;
wire n_0_0_110;
wire n_0_0_111;
wire n_0_0_112;
wire n_0_0_113;
wire n_0_0_114;
wire n_0_0_115;
wire n_0_0_116;
wire n_0_0_117;
wire n_0_0_118;
wire n_0_0_119;
wire n_0_0_120;
wire n_0_0_121;
wire n_0_0_122;
wire n_0_0_123;
wire n_0_0_124;
wire n_0_0_125;
wire n_0_0_126;
wire n_0_0_127;
wire n_0_0_128;
wire n_0_0_129;
wire n_0_0_130;
wire n_0_0_131;
wire n_0_0_132;
wire n_0_0_133;
wire n_0_0_134;
wire n_0_0_135;
wire n_0_0_136;
wire n_0_0_137;
wire n_0_0_138;
wire n_0_0_139;
wire n_0_0_140;
wire n_0_0_141;
wire n_0_0_142;
wire n_0_0_143;
wire n_0_0_144;
wire n_0_0_145;
wire n_0_0_146;
wire n_0_0_147;
wire n_0_0_148;
wire n_0_0_149;
wire n_0_0_150;
wire n_0_0_151;
wire n_0_0_152;
wire n_0_0_153;
wire n_0_0_154;
wire n_0_0_155;
wire n_0_0_156;
wire n_0_0_157;
wire n_0_0_158;
wire n_0_0_159;
wire n_0_0_160;
wire n_0_0_161;
wire n_0_0_162;
wire n_0_0_163;
wire n_0_0_164;
wire n_0_0_165;
wire n_0_0_166;
wire n_0_0_167;
wire n_0_0_168;
wire n_0_0_169;
wire n_0_0_170;
wire n_0_0_171;
wire n_0_0_172;
wire n_0_0_173;
wire n_0_0_174;
wire n_0_0_175;
wire n_0_0_176;
wire n_0_0_177;
wire n_0_0_178;
wire n_0_0_179;
wire n_0_0_180;
wire n_0_0_181;
wire n_0_0_182;
wire n_0_0_183;
wire n_0_0_184;
wire n_0_0_185;
wire n_0_0_186;
wire n_0_0_187;
wire n_0_0_188;
wire n_0_0_189;
wire n_0_0_190;
wire n_0_0_191;
wire n_0_0_192;
wire n_0_0_193;
wire n_0_0_194;
wire n_0_0_195;
wire n_0_0_196;
wire n_0_0_197;
wire n_0_0_198;
wire n_0_0_199;
wire n_0_0_200;
wire n_0_0_201;
wire n_0_0_202;
wire n_0_0_203;
wire n_0_0_204;
wire n_0_0_205;
wire n_0_0_206;
wire n_0_0_207;
wire n_0_0_208;
wire n_0_0_209;
wire n_0_0_210;
wire n_0_0_211;
wire n_0_0_212;
wire n_0_0_213;
wire n_0_0_214;
wire n_0_0_215;
wire n_0_0_216;
wire n_0_0_217;
wire n_0_0_218;
wire n_0_0_219;
wire n_0_0_220;
wire n_0_0_221;
wire n_0_0_222;
wire n_0_0_223;
wire n_0_0_224;
wire n_0_0_225;
wire n_0_0_226;
wire n_0_0_227;
wire n_0_0_228;
wire n_0_0_229;
wire n_0_0_230;
wire n_0_0_231;
wire n_0_0_232;
wire n_0_0_233;
wire n_0_0_234;
wire n_0_0_235;
wire n_0_0_236;
wire n_0_0_237;
wire n_0_0_238;
wire n_0_0_239;
wire n_0_0_240;
wire n_0_0_241;
wire n_0_0_242;
wire n_0_0_243;
wire n_0_0_244;
wire n_0_0_245;
wire n_0_0_246;
wire n_0_0_247;
wire n_0_0_248;
wire n_0_0_249;
wire n_0_0_250;
wire n_0_0_251;
wire n_0_0_252;
wire n_0_0_253;
wire n_0_0_254;
wire n_0_0_255;
wire n_0_0_256;
wire n_0_0_257;
wire n_0_0_258;
wire n_0_0_259;
wire n_0_0_260;
wire n_0_0_261;
wire n_0_0_262;
wire n_0_0_263;
wire n_0_0_264;
wire n_0_0_265;
wire n_0_0_266;
wire n_0_0_267;
wire n_0_0_268;
wire n_0_0_269;
wire n_0_0_270;
wire n_0_0_271;
wire n_0_0_272;
wire n_0_0_273;
wire n_0_0_274;
wire n_0_0_275;
wire n_0_0_276;
wire n_0_0_277;
wire n_0_0_278;
wire n_0_0_279;
wire n_0_0_280;
wire n_0_0_281;
wire n_0_0_282;
wire n_0_0_283;
wire n_0_0_284;
wire n_0_0_285;
wire n_0_0_286;
wire n_0_0_287;
wire n_0_0_288;
wire n_0_0_289;
wire n_0_0_290;
wire n_0_0_291;
wire n_0_0_292;
wire n_0_0_293;
wire n_0_0_294;
wire n_0_0_295;
wire n_0_0_296;
wire n_0_0_297;
wire n_0_0_298;
wire n_0_0_299;
wire n_0_0_300;
wire n_0_0_301;
wire n_0_0_302;
wire n_0_0_303;
wire n_0_0_304;
wire n_0_0_305;
wire n_0_0_306;
wire n_0_0_307;
wire n_0_0_308;
wire n_0_0_309;
wire n_0_0_310;
wire n_0_0_311;
wire n_0_0_312;
wire n_0_0_313;
wire n_0_0_314;
wire n_0_0_315;
wire n_0_0_316;
wire n_0_0_317;
wire n_0_0_318;
wire n_0_0_319;
wire n_0_0_320;
wire n_0_0_321;
wire n_0_0_322;
wire n_0_0_323;
wire n_0_0_324;
wire n_0_0_325;
wire n_0_0_326;
wire n_0_0_327;
wire n_0_0_328;
wire n_0_0_329;
wire n_0_0_330;
wire n_0_0_331;
wire n_0_0_332;
wire n_0_0_333;
wire n_0_0_334;
wire n_0_0_335;
wire n_0_0_336;
wire n_0_0_337;
wire n_0_0_338;
wire n_0_0_339;
wire n_0_0_340;
wire n_0_0_341;
wire n_0_0_342;
wire n_0_0_343;
wire n_0_0_344;
wire n_0_0_345;
wire n_0_0_346;
wire n_0_0_347;
wire n_0_0_348;
wire n_0_0_349;
wire n_0_0_350;
wire n_0_0_351;
wire n_0_0_352;
wire n_0_0_353;
wire n_0_0_354;
wire n_0_0_355;
wire n_0_0_356;
wire n_0_0_357;
wire n_0_0_358;
wire n_0_0_359;
wire n_0_0_360;
wire n_0_0_361;
wire n_0_0_362;
wire n_0_0_363;
wire n_0_0_364;
wire n_0_0_365;
wire n_0_0_366;
wire n_0_0_367;
wire n_0_0_368;
wire n_0_0_369;
wire n_0_0_370;
wire n_0_0_371;
wire n_0_0_372;
wire n_0_0_373;
wire n_0_0_374;
wire n_0_0_375;
wire n_0_0_376;
wire n_0_0_377;
wire n_0_0_378;
wire n_0_0_379;
wire n_0_0_380;
wire n_0_0_381;
wire n_0_0_382;
wire n_0_0_383;
wire n_0_0_384;
wire n_0_0_385;
wire n_0_0_386;
wire n_0_0_387;
wire n_0_0_388;
wire n_0_0_389;
wire n_0_0_390;
wire n_0_0_391;
wire n_0_0_392;
wire n_0_0_393;
wire n_0_0_394;
wire n_0_0_395;
wire n_0_0_396;
wire n_0_0_397;
wire n_0_0_398;
wire n_0_0_399;
wire n_0_0_400;
wire n_0_0_401;
wire n_0_0_402;
wire n_0_0_403;
wire n_0_0_404;
wire n_0_0_405;
wire n_0_0_406;
wire n_0_0_407;
wire n_0_0_408;
wire n_0_0_409;
wire n_0_0_410;
wire n_0_0_411;
wire n_0_0_412;
wire n_0_0_413;
wire n_0_0_414;
wire n_0_0_415;
wire n_0_0_416;
wire n_0_0_417;
wire n_0_0_418;
wire n_0_0_419;
wire n_0_0_420;
wire n_0_0_421;
wire n_0_0_422;
wire n_0_0_423;
wire n_0_0_424;
wire n_0_0_425;
wire n_0_0_426;
wire n_0_0_427;
wire n_0_0_428;
wire n_0_0_429;
wire n_0_0_430;
wire n_0_0_431;
wire n_0_0_432;
wire n_0_0_433;
wire n_0_0_434;
wire n_0_0_435;
wire n_0_0_436;
wire n_0_0_437;
wire n_0_0_438;
wire n_0_0_439;
wire n_0_0_440;
wire n_0_0_441;
wire n_0_0_442;
wire n_0_0_443;
wire n_0_0_444;
wire n_0_0_445;
wire n_0_0_446;
wire n_0_0_447;
wire n_0_0_448;
wire n_0_0_449;
wire n_0_0_450;
wire n_0_0_451;
wire n_0_0_452;
wire n_0_0_453;
wire n_0_0_454;
wire n_0_0_455;
wire n_0_0_456;
wire n_0_0_457;
wire n_0_0_458;
wire n_0_0_459;
wire n_0_0_460;
wire n_0_0_461;
wire n_0_0_462;
wire n_0_0_463;
wire n_0_0_464;
wire n_0_0_465;
wire n_0_0_466;
wire n_0_0_467;
wire n_0_0_468;
wire n_0_0_469;
wire n_0_0_470;
wire n_0_0_471;
wire n_0_0_472;
wire n_0_0_473;
wire n_0_0_474;
wire n_0_0_475;
wire n_0_0_476;
wire n_0_0_477;
wire n_0_0_478;
wire n_0_0_479;
wire n_0_0_480;
wire n_0_0_481;
wire n_0_0_482;
wire n_0_0_483;
wire n_0_0_484;
wire n_0_0_485;
wire n_0_0_486;
wire n_0_0_487;
wire n_0_0_488;
wire n_0_0_489;
wire n_0_0_490;
wire n_0_0_491;
wire n_0_0_492;
wire n_0_0_493;
wire n_0_0_494;
wire n_0_0_495;
wire n_0_0_496;
wire n_0_0_497;
wire n_0_0_498;
wire n_0_0_499;
wire n_0_0_500;
wire n_0_0_501;
wire n_0_0_502;
wire n_0_0_503;
wire n_0_0_504;
wire n_0_0_505;
wire n_0_0_506;
wire n_0_0_507;
wire n_0_0_508;
wire n_0_0_509;
wire n_0_0_510;
wire n_0_0_511;
wire n_0_0_512;
wire n_0_0_513;
wire n_0_0_514;
wire n_0_0_515;
wire n_0_0_516;
wire n_0_0_517;
wire n_0_0_518;
wire n_0_0_519;
wire n_0_0_520;
wire n_0_0_521;
wire n_0_0_522;
wire n_0_0_523;
wire n_0_0_524;
wire n_0_0_525;
wire n_0_0_526;
wire n_0_0_527;
wire n_0_0_528;
wire n_0_0_529;
wire n_0_0_530;
wire n_0_0_531;
wire n_0_0_532;
wire n_0_0_533;
wire n_0_0_534;
wire n_0_0_535;
wire n_0_0_536;
wire n_0_0_537;
wire n_0_0_538;
wire n_0_0_539;
wire n_0_0_540;
wire n_0_0_541;
wire n_0_0_542;
wire n_0_0_543;
wire n_0_0_544;
wire n_0_0_545;
wire n_0_0_546;
wire n_0_0_547;
wire n_0_0_548;
wire n_0_0_549;
wire n_0_0_550;
wire n_0_0_551;
wire n_0_0_552;
wire n_0_0_553;
wire n_0_0_554;
wire n_0_0_555;
wire n_0_0_556;
wire n_0_0_557;
wire n_0_0_558;
wire n_0_0_559;
wire n_0_0_560;
wire n_0_0_561;
wire n_0_0_562;
wire n_0_0_563;
wire n_0_0_564;
wire n_0_0_565;
wire n_0_0_566;
wire n_0_0_567;
wire n_0_0_568;
wire n_0_0_569;
wire n_0_0_570;
wire n_0_0_571;
wire n_0_0_572;
wire n_0_0_573;
wire n_0_0_574;
wire n_0_0_575;
wire n_0_0_576;
wire n_0_0_577;
wire n_0_0_578;
wire n_0_0_579;
wire n_0_0_580;
wire n_0_0_581;
wire n_0_0_582;
wire n_0_0_583;
wire n_0_0_584;
wire n_0_0_585;
wire n_0_0_586;
wire n_0_0_587;
wire n_0_0_588;
wire n_0_0_589;
wire n_0_0_590;
wire n_0_0_591;
wire n_0_0_592;
wire n_0_0_593;
wire n_0_0_594;
wire n_0_0_595;
wire n_0_0_596;
wire n_0_0_597;
wire n_0_0_598;
wire n_0_0_599;
wire n_0_0_600;
wire n_0_0_601;
wire n_0_0_602;
wire n_0_0_603;
wire n_0_0_604;
wire n_0_0_605;
wire n_0_0_606;
wire n_0_0_607;
wire n_0_0_608;
wire n_0_0_609;
wire n_0_0_610;
wire n_0_0_611;
wire n_0_0_612;
wire n_0_0_613;
wire n_0_0_614;
wire n_0_0_615;
wire n_0_0_616;
wire n_0_0_617;
wire n_0_0_618;
wire n_0_0_619;
wire n_0_0_620;
wire n_0_0_621;
wire n_0_0_622;
wire n_0_0_623;
wire n_0_0_624;
wire n_0_0_625;
wire n_0_0_626;
wire n_0_0_627;
wire n_0_0_628;
wire n_0_0_629;
wire n_0_0_630;
wire n_0_0_631;
wire n_0_0_632;
wire n_0_0_633;
wire n_0_0_634;
wire n_0_0_635;
wire n_0_0_636;
wire n_0_0_637;
wire n_0_0_638;
wire n_0_0_639;
wire n_0_0_640;
wire n_0_0_641;
wire n_0_0_642;
wire n_0_0_643;
wire n_0_0_644;
wire n_0_0_645;
wire n_0_0_646;
wire n_0_0_647;
wire n_0_0_648;
wire n_0_0_649;
wire n_0_0_650;
wire n_0_0_651;
wire n_0_0_652;
wire n_0_0_653;
wire n_0_0_654;
wire n_0_0_655;
wire n_0_0_656;
wire n_0_0_657;
wire n_0_0_658;
wire n_0_0_659;
wire n_0_0_660;
wire n_0_0_661;
wire n_0_0_662;
wire n_0_0_663;
wire n_0_0_664;
wire n_0_0_665;
wire n_0_0_666;
wire n_0_0_667;
wire n_0_0_668;
wire n_0_0_669;
wire n_0_0_670;
wire n_0_0_671;
wire n_0_0_672;
wire n_0_0_673;
wire n_0_0_674;
wire n_0_0_675;
wire n_0_0_676;
wire n_0_0_677;
wire n_0_0_678;
wire n_0_0_679;
wire n_0_0_680;
wire n_0_0_681;
wire n_0_0_682;
wire n_0_0_683;
wire n_0_0_684;
wire n_0_0_685;
wire n_0_0_686;
wire n_0_0_687;
wire n_0_0_688;
wire n_0_0_689;
wire n_0_0_690;
wire n_0_0_691;
wire n_0_0_692;
wire n_0_0_693;
wire n_0_0_694;
wire n_0_0_695;
wire n_0_0_696;
wire n_0_0_697;
wire n_0_0_698;
wire n_0_0_699;
wire n_0_0_700;
wire n_0_0_701;
wire n_0_0_702;
wire n_0_0_703;
wire n_0_0_704;
wire n_0_0_705;
wire n_0_0_706;
wire n_0_0_707;
wire n_0_0_708;
wire n_0_0_709;
wire n_0_0_710;
wire n_0_0_711;
wire n_0_0_712;
wire n_0_0_713;
wire n_0_0_714;
wire n_0_0_715;
wire n_0_0_716;
wire n_0_0_717;
wire n_0_0_718;
wire n_0_0_719;
wire n_0_0_720;
wire n_0_0_721;
wire n_0_0_722;
wire n_0_0_723;
wire n_0_0_724;
wire n_0_0_725;
wire n_0_0_726;
wire n_0_0_727;
wire n_0_0_728;
wire n_0_0_729;
wire n_0_0_730;
wire n_0_0_731;
wire n_0_0_732;
wire n_0_0_733;
wire n_0_0_734;
wire n_0_0_735;
wire n_0_0_736;
wire n_0_0_737;
wire n_0_0_738;
wire n_0_0_739;
wire n_0_0_740;
wire n_0_0_741;
wire n_0_0_742;
wire n_0_0_743;
wire n_0_0_744;
wire n_0_0_745;
wire n_0_0_746;
wire n_0_0_747;
wire n_0_0_748;
wire n_0_0_749;
wire n_0_0_750;
wire n_0_0_751;
wire n_0_0_752;
wire n_0_0_753;
wire n_0_0_754;
wire n_0_0_755;
wire n_0_0_756;
wire n_0_0_757;
wire n_0_0_758;
wire n_0_0_759;
wire n_0_0_760;
wire n_0_0_761;
wire n_0_0_762;
wire n_0_0_763;
wire n_0_0_764;
wire n_0_0_765;
wire n_0_0_766;
wire n_0_0_767;
wire n_0_0_768;
wire n_0_0_769;
wire n_0_0_770;
wire n_0_0_771;
wire n_0_0_772;
wire n_0_0_773;
wire n_0_0_774;
wire n_0_0_775;
wire n_0_0_776;
wire n_0_0_777;
wire n_0_0_778;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_0_779;
wire n_0_164;
wire n_0_160;
wire n_0_165;
wire n_0_166;
wire \Acc[63] ;
wire \Acc[62] ;
wire \Acc[61] ;
wire \Acc[60] ;
wire \Acc[59] ;
wire \Acc[58] ;
wire \Acc[57] ;
wire \Acc[56] ;
wire \Acc[55] ;
wire \Acc[54] ;
wire \Acc[53] ;
wire \Acc[52] ;
wire \Acc[51] ;
wire \Acc[50] ;
wire \Acc[49] ;
wire \Acc[48] ;
wire \Acc[47] ;
wire \Acc[46] ;
wire \Acc[45] ;
wire \Acc[44] ;
wire \Acc[43] ;
wire \Acc[42] ;
wire \Acc[41] ;
wire \Acc[40] ;
wire \Acc[39] ;
wire \Acc[38] ;
wire \Acc[37] ;
wire \Acc[36] ;
wire \Acc[35] ;
wire \Acc[34] ;
wire \Acc[33] ;
wire \Acc[32] ;
wire \Acc[31] ;
wire \Acc[30] ;
wire \Acc[29] ;
wire \Acc[28] ;
wire \Acc[27] ;
wire \Acc[26] ;
wire \Acc[25] ;
wire \Acc[24] ;
wire \Acc[23] ;
wire \Acc[22] ;
wire \Acc[21] ;
wire \Acc[20] ;
wire \Acc[19] ;
wire \Acc[18] ;
wire \Acc[17] ;
wire \Acc[16] ;
wire \Acc[15] ;
wire \Acc[14] ;
wire \Acc[13] ;
wire \Acc[12] ;
wire \Acc[11] ;
wire \Acc[10] ;
wire \Acc[9] ;
wire \Acc[8] ;
wire \Acc[7] ;
wire \Acc[6] ;
wire \Acc[5] ;
wire \Acc[4] ;
wire \Acc[3] ;
wire \Acc[2] ;
wire \Acc[1] ;
wire \Acc[0] ;
wire \i[5] ;
wire \i[4] ;
wire \i[3] ;
wire \i[2] ;
wire \i[1] ;
wire \Q[32] ;
wire \Q[31] ;
wire \Q[30] ;
wire \Q[29] ;
wire \Q[28] ;
wire \Q[27] ;
wire \Q[26] ;
wire \Q[25] ;
wire \Q[24] ;
wire \Q[23] ;
wire \Q[22] ;
wire \Q[21] ;
wire \Q[20] ;
wire \Q[19] ;
wire \Q[18] ;
wire \Q[17] ;
wire \Q[16] ;
wire \Q[15] ;
wire \Q[14] ;
wire \Q[13] ;
wire \Q[12] ;
wire \Q[11] ;
wire \Q[10] ;
wire \Q[9] ;
wire \Q[8] ;
wire \Q[7] ;
wire \Q[6] ;
wire \Q[5] ;
wire \Q[4] ;
wire \Q[3] ;
wire \Q[2] ;
wire \Q[1] ;
wire CTS_n98;
wire \extended_M_mul_neg_one[63] ;
wire CTS_n188;
wire CTS_n190;
wire \extended_M_mul_neg_one[30] ;
wire \extended_M_mul_neg_one[29] ;
wire \extended_M_mul_neg_one[28] ;
wire \extended_M_mul_neg_one[27] ;
wire \extended_M_mul_neg_one[26] ;
wire \extended_M_mul_neg_one[25] ;
wire \extended_M_mul_neg_one[24] ;
wire \extended_M_mul_neg_one[23] ;
wire \extended_M_mul_neg_one[22] ;
wire \extended_M_mul_neg_one[21] ;
wire \extended_M_mul_neg_one[20] ;
wire \extended_M_mul_neg_one[19] ;
wire \extended_M_mul_neg_one[18] ;
wire \extended_M_mul_neg_one[17] ;
wire \extended_M_mul_neg_one[16] ;
wire \extended_M_mul_neg_one[15] ;
wire \extended_M_mul_neg_one[14] ;
wire \extended_M_mul_neg_one[13] ;
wire \extended_M_mul_neg_one[12] ;
wire \extended_M_mul_neg_one[11] ;
wire \extended_M_mul_neg_one[10] ;
wire \extended_M_mul_neg_one[9] ;
wire \extended_M_mul_neg_one[8] ;
wire \extended_M_mul_neg_one[7] ;
wire \extended_M_mul_neg_one[6] ;
wire \extended_M_mul_neg_one[5] ;
wire \extended_M_mul_neg_one[4] ;
wire \extended_M_mul_neg_one[3] ;
wire \extended_M_mul_neg_one[2] ;
wire \extended_M_mul_neg_one[1] ;
wire CTS_n189;
wire \extended_M[63] ;
wire CLOCK_n311;
wire CTS_n215;
wire hfn_ipo_n67;
wire drc_ipo_n84;
wire hfn_ipo_n80;
wire hfn_ipo_n79;
wire hfn_ipo_n78;
wire hfn_ipo_n77;
wire hfn_ipo_n73;
wire CTS_n146;
wire hfn_ipo_n69;
wire hfn_ipo_n71;
wire CTS_n187;
wire hfn_ipo_n64;
wire hfn_ipo_n63;
wire hfn_ipo_n62;
wire hfn_ipo_n61;
wire hfn_ipo_n66;
wire hfn_ipo_n65;
wire hfn_ipo_n60;
wire hfn_ipo_n59;
wire drc_ipo_n83;
wire hfn_ipo_n82;
wire hfn_ipo_n81;
wire hfn_ipo_n76;
wire hfn_ipo_n75;
wire CTS_n285;
wire CTS_n99;
wire hfn_ipo_n57;
wire \extended_M[30] ;
wire \extended_M[29] ;
wire \extended_M[28] ;
wire \extended_M[27] ;
wire \extended_M[26] ;
wire \extended_M[25] ;
wire \extended_M[24] ;
wire \extended_M[23] ;
wire \extended_M[22] ;
wire \extended_M[21] ;
wire \extended_M[20] ;
wire \extended_M[19] ;
wire \extended_M[18] ;
wire \extended_M[17] ;
wire \extended_M[16] ;
wire \extended_M[15] ;
wire \extended_M[14] ;
wire \extended_M[13] ;
wire \extended_M[12] ;
wire \extended_M[11] ;
wire \extended_M[10] ;
wire \extended_M[9] ;
wire \extended_M[8] ;
wire \extended_M[7] ;
wire \extended_M[6] ;
wire \extended_M[5] ;
wire \extended_M[4] ;
wire \extended_M[3] ;
wire \extended_M[2] ;
wire \extended_M[1] ;
wire \extended_M[0] ;
wire uc_0;


DFF_X1 \extended_M_reg[63]  (.Q (\extended_M[63] ), .CK (CTS_n98), .D (\A_reg[31] ));
DFF_X1 \extended_M_mul_neg_one_reg[63]  (.Q (\extended_M_mul_neg_one[63] ), .CK (CTS_n98), .D (n_0_32));
DFF_X1 \extended_M_reg[0]  (.Q (\extended_M[0] ), .CK (CTS_n99), .D (\A_reg[0] ));
DFF_X1 \extended_M_reg[30]  (.Q (\extended_M[30] ), .CK (CTS_n98), .D (\A_reg[30] ));
DFF_X1 \extended_M_reg[14]  (.Q (\extended_M[14] ), .CK (CTS_n98), .D (\A_reg[14] ));
DFF_X1 \extended_M_reg[22]  (.Q (\extended_M[22] ), .CK (CTS_n99), .D (\A_reg[22] ));
DFF_X1 \extended_M_reg[6]  (.Q (\extended_M[6] ), .CK (CTS_n99), .D (\A_reg[6] ));
DFF_X1 \extended_M_reg[26]  (.Q (\extended_M[26] ), .CK (CTS_n98), .D (\A_reg[26] ));
DFF_X1 \extended_M_reg[10]  (.Q (\extended_M[10] ), .CK (CTS_n99), .D (\A_reg[10] ));
DFF_X1 \extended_M_reg[18]  (.Q (\extended_M[18] ), .CK (CTS_n99), .D (\A_reg[18] ));
DFF_X1 \extended_M_reg[2]  (.Q (\extended_M[2] ), .CK (CTS_n99), .D (\A_reg[2] ));
DFF_X1 \extended_M_reg[28]  (.Q (\extended_M[28] ), .CK (CTS_n98), .D (\A_reg[28] ));
DFF_X1 \extended_M_reg[12]  (.Q (\extended_M[12] ), .CK (CTS_n99), .D (\A_reg[12] ));
DFF_X1 \extended_M_reg[20]  (.Q (\extended_M[20] ), .CK (CTS_n99), .D (\A_reg[20] ));
DFF_X1 \extended_M_reg[4]  (.Q (\extended_M[4] ), .CK (CTS_n99), .D (\A_reg[4] ));
DFF_X1 \extended_M_reg[24]  (.Q (\extended_M[24] ), .CK (CTS_n99), .D (\A_reg[24] ));
DFF_X1 \extended_M_reg[8]  (.Q (\extended_M[8] ), .CK (CTS_n99), .D (\A_reg[8] ));
DFF_X1 \extended_M_reg[16]  (.Q (\extended_M[16] ), .CK (CTS_n99), .D (\A_reg[16] ));
DFF_X1 \extended_M_reg[29]  (.Q (\extended_M[29] ), .CK (CTS_n98), .D (\A_reg[29] ));
DFF_X1 \extended_M_reg[13]  (.Q (\extended_M[13] ), .CK (CTS_n99), .D (\A_reg[13] ));
DFF_X1 \extended_M_reg[21]  (.Q (\extended_M[21] ), .CK (CTS_n99), .D (\A_reg[21] ));
DFF_X1 \extended_M_reg[5]  (.Q (\extended_M[5] ), .CK (CTS_n99), .D (\A_reg[5] ));
DFF_X1 \extended_M_reg[25]  (.Q (\extended_M[25] ), .CK (CTS_n99), .D (\A_reg[25] ));
DFF_X1 \extended_M_reg[9]  (.Q (\extended_M[9] ), .CK (CTS_n99), .D (\A_reg[9] ));
DFF_X1 \extended_M_reg[17]  (.Q (\extended_M[17] ), .CK (CTS_n99), .D (\A_reg[17] ));
DFF_X1 \extended_M_reg[1]  (.Q (\extended_M[1] ), .CK (CTS_n99), .D (\A_reg[1] ));
DFF_X1 \extended_M_reg[27]  (.Q (\extended_M[27] ), .CK (CTS_n98), .D (\A_reg[27] ));
DFF_X1 \extended_M_reg[11]  (.Q (\extended_M[11] ), .CK (CTS_n99), .D (\A_reg[11] ));
DFF_X1 \extended_M_reg[19]  (.Q (\extended_M[19] ), .CK (CTS_n99), .D (\A_reg[19] ));
DFF_X1 \extended_M_reg[3]  (.Q (\extended_M[3] ), .CK (CTS_n99), .D (\A_reg[3] ));
DFF_X1 \extended_M_reg[23]  (.Q (\extended_M[23] ), .CK (CTS_n99), .D (\A_reg[23] ));
DFF_X1 \extended_M_reg[7]  (.Q (\extended_M[7] ), .CK (CTS_n99), .D (\A_reg[7] ));
DFF_X1 \extended_M_reg[15]  (.Q (\extended_M[15] ), .CK (CTS_n99), .D (\A_reg[15] ));
DFF_X1 \extended_M_mul_neg_one_reg[30]  (.Q (\extended_M_mul_neg_one[30] ), .CK (CTS_n98), .D (n_0_31));
DFF_X1 \extended_M_mul_neg_one_reg[14]  (.Q (\extended_M_mul_neg_one[14] ), .CK (CTS_n98), .D (n_0_15));
DFF_X1 \extended_M_mul_neg_one_reg[22]  (.Q (\extended_M_mul_neg_one[22] ), .CK (CTS_n99), .D (n_0_23));
DFF_X1 \extended_M_mul_neg_one_reg[6]  (.Q (\extended_M_mul_neg_one[6] ), .CK (CTS_n99), .D (n_0_7));
DFF_X1 \extended_M_mul_neg_one_reg[26]  (.Q (\extended_M_mul_neg_one[26] ), .CK (CTS_n98), .D (n_0_27));
DFF_X1 \extended_M_mul_neg_one_reg[10]  (.Q (\extended_M_mul_neg_one[10] ), .CK (CTS_n99), .D (n_0_11));
DFF_X1 \extended_M_mul_neg_one_reg[18]  (.Q (\extended_M_mul_neg_one[18] ), .CK (CTS_n99), .D (n_0_19));
DFF_X1 \extended_M_mul_neg_one_reg[2]  (.Q (\extended_M_mul_neg_one[2] ), .CK (CTS_n99), .D (n_0_3));
DFF_X1 \extended_M_mul_neg_one_reg[28]  (.Q (\extended_M_mul_neg_one[28] ), .CK (CTS_n98), .D (n_0_29));
DFF_X1 \extended_M_mul_neg_one_reg[12]  (.Q (\extended_M_mul_neg_one[12] ), .CK (CTS_n98), .D (n_0_13));
DFF_X1 \extended_M_mul_neg_one_reg[20]  (.Q (\extended_M_mul_neg_one[20] ), .CK (CTS_n99), .D (n_0_21));
DFF_X1 \extended_M_mul_neg_one_reg[4]  (.Q (\extended_M_mul_neg_one[4] ), .CK (CTS_n99), .D (n_0_5));
DFF_X1 \extended_M_mul_neg_one_reg[24]  (.Q (\extended_M_mul_neg_one[24] ), .CK (CTS_n99), .D (n_0_25));
DFF_X1 \extended_M_mul_neg_one_reg[8]  (.Q (\extended_M_mul_neg_one[8] ), .CK (CTS_n99), .D (n_0_9));
DFF_X1 \extended_M_mul_neg_one_reg[16]  (.Q (\extended_M_mul_neg_one[16] ), .CK (CTS_n99), .D (n_0_17));
DFF_X1 \extended_M_mul_neg_one_reg[29]  (.Q (\extended_M_mul_neg_one[29] ), .CK (CTS_n98), .D (n_0_30));
DFF_X1 \extended_M_mul_neg_one_reg[13]  (.Q (\extended_M_mul_neg_one[13] ), .CK (CTS_n98), .D (n_0_14));
DFF_X1 \extended_M_mul_neg_one_reg[21]  (.Q (\extended_M_mul_neg_one[21] ), .CK (CTS_n99), .D (n_0_22));
DFF_X1 \extended_M_mul_neg_one_reg[5]  (.Q (\extended_M_mul_neg_one[5] ), .CK (CTS_n99), .D (n_0_6));
DFF_X1 \extended_M_mul_neg_one_reg[25]  (.Q (\extended_M_mul_neg_one[25] ), .CK (CTS_n99), .D (n_0_26));
DFF_X1 \extended_M_mul_neg_one_reg[9]  (.Q (\extended_M_mul_neg_one[9] ), .CK (CTS_n99), .D (n_0_10));
DFF_X1 \extended_M_mul_neg_one_reg[17]  (.Q (\extended_M_mul_neg_one[17] ), .CK (CTS_n99), .D (n_0_18));
DFF_X1 \extended_M_mul_neg_one_reg[1]  (.Q (\extended_M_mul_neg_one[1] ), .CK (CTS_n99), .D (n_0_2));
DFF_X1 \extended_M_mul_neg_one_reg[27]  (.Q (\extended_M_mul_neg_one[27] ), .CK (CTS_n98), .D (n_0_28));
DFF_X1 \extended_M_mul_neg_one_reg[11]  (.Q (\extended_M_mul_neg_one[11] ), .CK (CTS_n99), .D (n_0_12));
DFF_X1 \extended_M_mul_neg_one_reg[19]  (.Q (\extended_M_mul_neg_one[19] ), .CK (CTS_n99), .D (n_0_20));
DFF_X1 \extended_M_mul_neg_one_reg[3]  (.Q (\extended_M_mul_neg_one[3] ), .CK (CTS_n99), .D (n_0_4));
DFF_X1 \extended_M_mul_neg_one_reg[23]  (.Q (\extended_M_mul_neg_one[23] ), .CK (CTS_n99), .D (n_0_24));
DFF_X1 \extended_M_mul_neg_one_reg[7]  (.Q (\extended_M_mul_neg_one[7] ), .CK (CTS_n99), .D (n_0_8));
DFF_X1 \extended_M_mul_neg_one_reg[15]  (.Q (\extended_M_mul_neg_one[15] ), .CK (CTS_n99), .D (n_0_16));
CLKGATETST_X8 clk_gate_extended_M_reg (.GCK (CTS_n146), .CK (CTS_n285), .E (start), .SE (VSS));
CLKGATETST_X4 clk_gate_Acc_reg (.GCK (CTS_n187), .CK (CLOCK_n311), .E (n_0_165), .SE (VSS));
DFF_X1 \Q_reg[1]  (.Q (\Q[1] ), .CK (CTS_n98), .D (\B_reg[0] ));
DFF_X1 \Q_reg[2]  (.Q (\Q[2] ), .CK (CTS_n98), .D (\B_reg[1] ));
DFF_X1 \Q_reg[3]  (.Q (\Q[3] ), .CK (CTS_n98), .D (\B_reg[2] ));
DFF_X1 \Q_reg[4]  (.Q (\Q[4] ), .CK (CTS_n98), .D (\B_reg[3] ));
DFF_X1 \Q_reg[5]  (.Q (\Q[5] ), .CK (CTS_n98), .D (\B_reg[4] ));
DFF_X1 \Q_reg[6]  (.Q (\Q[6] ), .CK (CTS_n98), .D (\B_reg[5] ));
DFF_X1 \Q_reg[7]  (.Q (\Q[7] ), .CK (CTS_n98), .D (\B_reg[6] ));
DFF_X1 \Q_reg[8]  (.Q (\Q[8] ), .CK (CTS_n98), .D (\B_reg[7] ));
DFF_X1 \Q_reg[9]  (.Q (\Q[9] ), .CK (CTS_n98), .D (\B_reg[8] ));
DFF_X1 \Q_reg[10]  (.Q (\Q[10] ), .CK (CTS_n98), .D (\B_reg[9] ));
DFF_X1 \Q_reg[11]  (.Q (\Q[11] ), .CK (CTS_n98), .D (\B_reg[10] ));
DFF_X1 \Q_reg[12]  (.Q (\Q[12] ), .CK (CTS_n98), .D (\B_reg[11] ));
DFF_X1 \Q_reg[13]  (.Q (\Q[13] ), .CK (CTS_n98), .D (\B_reg[12] ));
DFF_X1 \Q_reg[14]  (.Q (\Q[14] ), .CK (CTS_n98), .D (\B_reg[13] ));
DFF_X1 \Q_reg[15]  (.Q (\Q[15] ), .CK (CTS_n98), .D (\B_reg[14] ));
DFF_X1 \Q_reg[16]  (.Q (\Q[16] ), .CK (CTS_n98), .D (\B_reg[15] ));
DFF_X1 \Q_reg[17]  (.Q (\Q[17] ), .CK (CTS_n98), .D (\B_reg[16] ));
DFF_X1 \Q_reg[18]  (.Q (\Q[18] ), .CK (CTS_n98), .D (\B_reg[17] ));
DFF_X1 \Q_reg[19]  (.Q (\Q[19] ), .CK (CTS_n98), .D (\B_reg[18] ));
DFF_X1 \Q_reg[20]  (.Q (\Q[20] ), .CK (CTS_n98), .D (\B_reg[19] ));
DFF_X1 \Q_reg[21]  (.Q (\Q[21] ), .CK (CTS_n98), .D (\B_reg[20] ));
DFF_X1 \Q_reg[22]  (.Q (\Q[22] ), .CK (CTS_n98), .D (\B_reg[21] ));
DFF_X1 \Q_reg[23]  (.Q (\Q[23] ), .CK (CTS_n98), .D (\B_reg[22] ));
DFF_X1 \Q_reg[24]  (.Q (\Q[24] ), .CK (CTS_n98), .D (\B_reg[23] ));
DFF_X1 \Q_reg[25]  (.Q (\Q[25] ), .CK (CTS_n98), .D (\B_reg[24] ));
DFF_X1 \Q_reg[26]  (.Q (\Q[26] ), .CK (CTS_n98), .D (\B_reg[25] ));
DFF_X1 \Q_reg[27]  (.Q (\Q[27] ), .CK (CTS_n98), .D (\B_reg[26] ));
DFF_X1 \Q_reg[28]  (.Q (\Q[28] ), .CK (CTS_n98), .D (\B_reg[27] ));
DFF_X1 \Q_reg[29]  (.Q (\Q[29] ), .CK (CTS_n98), .D (\B_reg[28] ));
DFF_X1 \Q_reg[30]  (.Q (\Q[30] ), .CK (CTS_n98), .D (\B_reg[29] ));
DFF_X1 \Q_reg[31]  (.Q (\Q[31] ), .CK (CTS_n98), .D (\B_reg[30] ));
DFF_X1 \Q_reg[32]  (.Q (\Q[32] ), .CK (CTS_n98), .D (\B_reg[31] ));
DFF_X1 \i_reg[1]  (.Q (\i[1] ), .CK (CTS_n189), .D (n_0_160));
DFF_X1 \i_reg[2]  (.Q (\i[2] ), .CK (CTS_n189), .D (n_0_161));
DFF_X1 \i_reg[3]  (.Q (\i[3] ), .CK (CTS_n189), .D (n_0_162));
DFF_X1 \i_reg[4]  (.Q (\i[4] ), .CK (CTS_n189), .D (n_0_163));
DFF_X1 \i_reg[5]  (.Q (\i[5] ), .CK (CTS_n189), .D (n_0_164));
DFF_X1 \Acc_reg[0]  (.Q (\Acc[0] ), .CK (CTS_n189), .D (n_0_96));
DFF_X1 \Acc_reg[1]  (.Q (\Acc[1] ), .CK (CTS_n189), .D (n_0_97));
DFF_X1 \Acc_reg[2]  (.Q (\Acc[2] ), .CK (CTS_n189), .D (n_0_98));
DFF_X1 \Acc_reg[3]  (.Q (\Acc[3] ), .CK (CTS_n189), .D (n_0_99));
DFF_X1 \Acc_reg[4]  (.Q (\Acc[4] ), .CK (CTS_n189), .D (n_0_100));
DFF_X1 \Acc_reg[5]  (.Q (\Acc[5] ), .CK (CTS_n189), .D (n_0_101));
DFF_X1 \Acc_reg[6]  (.Q (\Acc[6] ), .CK (CTS_n189), .D (n_0_102));
DFF_X1 \Acc_reg[7]  (.Q (\Acc[7] ), .CK (CTS_n189), .D (n_0_103));
DFF_X1 \Acc_reg[8]  (.Q (\Acc[8] ), .CK (CTS_n189), .D (n_0_104));
DFF_X1 \Acc_reg[9]  (.Q (\Acc[9] ), .CK (CTS_n189), .D (n_0_105));
DFF_X1 \Acc_reg[10]  (.Q (\Acc[10] ), .CK (CTS_n189), .D (n_0_106));
DFF_X1 \Acc_reg[11]  (.Q (\Acc[11] ), .CK (CTS_n189), .D (n_0_107));
DFF_X1 \Acc_reg[12]  (.Q (\Acc[12] ), .CK (CTS_n189), .D (n_0_108));
DFF_X1 \Acc_reg[13]  (.Q (\Acc[13] ), .CK (CTS_n189), .D (n_0_109));
DFF_X1 \Acc_reg[14]  (.Q (\Acc[14] ), .CK (CTS_n189), .D (n_0_110));
DFF_X1 \Acc_reg[15]  (.Q (\Acc[15] ), .CK (CTS_n189), .D (n_0_111));
DFF_X1 \Acc_reg[16]  (.Q (\Acc[16] ), .CK (CTS_n189), .D (n_0_112));
DFF_X1 \Acc_reg[17]  (.Q (\Acc[17] ), .CK (CTS_n189), .D (n_0_113));
DFF_X1 \Acc_reg[18]  (.Q (\Acc[18] ), .CK (CTS_n189), .D (n_0_114));
DFF_X1 \Acc_reg[19]  (.Q (\Acc[19] ), .CK (CTS_n190), .D (n_0_115));
DFF_X1 \Acc_reg[20]  (.Q (\Acc[20] ), .CK (CTS_n190), .D (n_0_116));
DFF_X1 \Acc_reg[21]  (.Q (\Acc[21] ), .CK (CTS_n190), .D (n_0_117));
DFF_X1 \Acc_reg[22]  (.Q (\Acc[22] ), .CK (CTS_n190), .D (n_0_118));
DFF_X1 \Acc_reg[23]  (.Q (\Acc[23] ), .CK (CTS_n190), .D (n_0_119));
DFF_X1 \Acc_reg[24]  (.Q (\Acc[24] ), .CK (CTS_n190), .D (n_0_120));
DFF_X1 \Acc_reg[25]  (.Q (\Acc[25] ), .CK (CTS_n190), .D (n_0_121));
DFF_X1 \Acc_reg[26]  (.Q (\Acc[26] ), .CK (CTS_n190), .D (n_0_122));
DFF_X1 \Acc_reg[27]  (.Q (\Acc[27] ), .CK (CTS_n190), .D (n_0_123));
DFF_X1 \Acc_reg[28]  (.Q (\Acc[28] ), .CK (CTS_n190), .D (n_0_124));
DFF_X1 \Acc_reg[29]  (.Q (\Acc[29] ), .CK (CTS_n190), .D (n_0_125));
DFF_X1 \Acc_reg[30]  (.Q (\Acc[30] ), .CK (CTS_n190), .D (n_0_126));
DFF_X1 \Acc_reg[31]  (.Q (\Acc[31] ), .CK (CTS_n190), .D (n_0_127));
DFF_X1 \Acc_reg[32]  (.Q (\Acc[32] ), .CK (CTS_n190), .D (n_0_128));
DFF_X1 \Acc_reg[33]  (.Q (\Acc[33] ), .CK (CTS_n190), .D (n_0_129));
DFF_X1 \Acc_reg[34]  (.Q (\Acc[34] ), .CK (CTS_n190), .D (n_0_130));
DFF_X1 \Acc_reg[35]  (.Q (\Acc[35] ), .CK (CTS_n190), .D (n_0_131));
DFF_X1 \Acc_reg[36]  (.Q (\Acc[36] ), .CK (CTS_n190), .D (n_0_132));
DFF_X1 \Acc_reg[37]  (.Q (\Acc[37] ), .CK (CTS_n190), .D (n_0_133));
DFF_X1 \Acc_reg[38]  (.Q (\Acc[38] ), .CK (CTS_n190), .D (n_0_134));
DFF_X1 \Acc_reg[39]  (.Q (\Acc[39] ), .CK (CTS_n190), .D (n_0_135));
DFF_X1 \Acc_reg[40]  (.Q (\Acc[40] ), .CK (CTS_n190), .D (n_0_136));
DFF_X1 \Acc_reg[41]  (.Q (\Acc[41] ), .CK (CTS_n188), .D (n_0_137));
DFF_X1 \Acc_reg[42]  (.Q (\Acc[42] ), .CK (CTS_n188), .D (n_0_138));
DFF_X1 \Acc_reg[43]  (.Q (\Acc[43] ), .CK (CTS_n188), .D (n_0_139));
DFF_X1 \Acc_reg[44]  (.Q (\Acc[44] ), .CK (CTS_n188), .D (n_0_140));
DFF_X1 \Acc_reg[45]  (.Q (\Acc[45] ), .CK (CTS_n188), .D (n_0_141));
DFF_X1 \Acc_reg[46]  (.Q (\Acc[46] ), .CK (CTS_n188), .D (n_0_142));
DFF_X1 \Acc_reg[47]  (.Q (\Acc[47] ), .CK (CTS_n188), .D (n_0_143));
DFF_X1 \Acc_reg[48]  (.Q (\Acc[48] ), .CK (CTS_n188), .D (n_0_144));
DFF_X1 \Acc_reg[49]  (.Q (\Acc[49] ), .CK (CTS_n188), .D (n_0_145));
DFF_X1 \Acc_reg[50]  (.Q (\Acc[50] ), .CK (CTS_n189), .D (n_0_146));
DFF_X1 \Acc_reg[51]  (.Q (\Acc[51] ), .CK (CTS_n189), .D (n_0_147));
DFF_X1 \Acc_reg[52]  (.Q (\Acc[52] ), .CK (CTS_n189), .D (n_0_148));
DFF_X1 \Acc_reg[53]  (.Q (\Acc[53] ), .CK (CTS_n189), .D (n_0_149));
DFF_X1 \Acc_reg[54]  (.Q (\Acc[54] ), .CK (CTS_n188), .D (n_0_150));
DFF_X1 \Acc_reg[55]  (.Q (\Acc[55] ), .CK (CTS_n188), .D (n_0_151));
DFF_X1 \Acc_reg[56]  (.Q (\Acc[56] ), .CK (CTS_n188), .D (n_0_152));
DFF_X1 \Acc_reg[57]  (.Q (\Acc[57] ), .CK (CTS_n188), .D (n_0_153));
DFF_X1 \Acc_reg[58]  (.Q (\Acc[58] ), .CK (CTS_n188), .D (n_0_154));
DFF_X1 \Acc_reg[59]  (.Q (\Acc[59] ), .CK (CTS_n188), .D (n_0_155));
DFF_X1 \Acc_reg[60]  (.Q (\Acc[60] ), .CK (CTS_n188), .D (n_0_156));
DFF_X1 \Acc_reg[61]  (.Q (\Acc[61] ), .CK (CTS_n188), .D (n_0_157));
DFF_X1 \Acc_reg[62]  (.Q (\Acc[62] ), .CK (CTS_n188), .D (n_0_158));
DFF_X1 \Acc_reg[63]  (.Q (\Acc[63] ), .CK (CTS_n188), .D (n_0_159));
INV_X1 i_0_0_911 (.ZN (n_0_166), .A (n_0_165));
NAND3_X1 i_0_0_910 (.ZN (n_0_165), .A1 (n_0_0_47), .A2 (n_0_0_20), .A3 (n_0_160));
NOR2_X1 i_0_0_909 (.ZN (n_0_160), .A1 (CLOCK_slh_n317), .A2 (hfn_ipo_n80));
AOI221_X1 i_0_0_908 (.ZN (n_0_164), .A (CLOCK_slh_n317), .B1 (drc_ipo_n84), .B2 (n_0_0_2)
    , .C1 (n_0_0_7), .C2 (n_0_0_779));
INV_X1 i_0_0_907 (.ZN (n_0_0_779), .A (n_0_0_2));
AND2_X1 i_0_0_906 (.ZN (n_0_163), .A1 (n_0_0_6), .A2 (n_0_0_5));
AND2_X1 i_0_0_905 (.ZN (n_0_162), .A1 (n_0_0_6), .A2 (n_0_0_4));
AND2_X1 i_0_0_904 (.ZN (n_0_161), .A1 (n_0_0_6), .A2 (n_0_0_3));
OAI21_X1 i_0_0_903 (.ZN (\partialProd[63] ), .A (n_0_0_765), .B1 (n_0_0_73), .B2 (n_0_0_778));
OAI21_X1 i_0_0_902 (.ZN (n_0_0_778), .A (n_0_0_777), .B1 (n_0_0_761), .B2 (hfn_ipo_n62));
OAI221_X1 i_0_0_901 (.ZN (n_0_0_777), .A (hfn_ipo_n63), .B1 (n_0_0_775), .B2 (n_0_0_776)
    , .C1 (n_0_0_737), .C2 (hfn_ipo_n59));
AOI21_X1 i_0_0_900 (.ZN (n_0_0_776), .A (hfn_ipo_n73), .B1 (n_0_0_694), .B2 (n_0_0_766));
OAI21_X1 i_0_0_899 (.ZN (n_0_0_775), .A (hfn_ipo_n59), .B1 (n_0_0_774), .B2 (hfn_ipo_n75));
OAI22_X1 i_0_0_898 (.ZN (n_0_0_774), .A1 (n_0_0_773), .A2 (n_0_0_664), .B1 (n_0_0_772), .B2 (n_0_0_213));
INV_X1 i_0_0_897 (.ZN (n_0_0_773), .A (n_0_0_772));
NAND2_X1 i_0_0_896 (.ZN (n_0_0_772), .A1 (drc_ipo_n83), .A2 (drc_ipo_n84));
OAI21_X1 i_0_0_895 (.ZN (\partialProd[62] ), .A (n_0_0_765), .B1 (n_0_0_73), .B2 (n_0_0_771));
OAI21_X1 i_0_0_894 (.ZN (n_0_0_771), .A (n_0_0_769), .B1 (n_0_0_770), .B2 (hfn_ipo_n62));
INV_X1 i_0_0_893 (.ZN (n_0_0_770), .A (n_0_0_751));
OAI211_X1 i_0_0_892 (.ZN (n_0_0_769), .A (hfn_ipo_n62), .B (n_0_0_767), .C1 (n_0_0_768), .C2 (hfn_ipo_n59));
INV_X1 i_0_0_891 (.ZN (n_0_0_768), .A (n_0_0_728));
OAI211_X1 i_0_0_890 (.ZN (n_0_0_767), .A (hfn_ipo_n59), .B (n_0_0_766), .C1 (n_0_0_420), .C2 (n_0_0_7));
INV_X1 i_0_0_889 (.ZN (n_0_0_766), .A (n_0_0_460));
AOI221_X1 i_0_0_888 (.ZN (n_0_0_765), .A (n_0_0_758), .B1 (hfn_ipo_n71), .B2 (n_0_0_763)
    , .C1 (hfn_ipo_n69), .C2 (n_0_0_757));
NAND2_X1 i_0_0_887 (.ZN (\partialProd[61] ), .A1 (n_0_0_759), .A2 (n_0_0_764));
AOI22_X1 i_0_0_886 (.ZN (n_0_0_764), .A1 (hfn_ipo_n67), .A2 (n_0_0_763), .B1 (hfn_ipo_n69), .B2 (n_0_0_748));
AOI22_X1 i_0_0_885 (.ZN (n_0_0_763), .A1 (n_0_0_739), .A2 (hfn_ipo_n80), .B1 (n_0_0_762), .B2 (hfn_ipo_n62));
INV_X1 i_0_0_884 (.ZN (n_0_0_762), .A (n_0_0_761));
AOI21_X1 i_0_0_883 (.ZN (n_0_0_761), .A (n_0_0_760), .B1 (hfn_ipo_n78), .B2 (n_0_0_722));
AOI211_X1 i_0_0_882 (.ZN (n_0_0_760), .A (hfn_ipo_n78), .B (n_0_0_614), .C1 (n_0_0_406), .C2 (drc_ipo_n84));
AOI21_X1 i_0_0_881 (.ZN (n_0_0_759), .A (n_0_0_758), .B1 (hfn_ipo_n71), .B2 (n_0_0_752));
AND2_X1 i_0_0_880 (.ZN (n_0_0_758), .A1 (hfn_ipo_n65), .A2 (n_0_0_757));
OAI22_X1 i_0_0_879 (.ZN (n_0_0_757), .A1 (n_0_0_756), .A2 (hfn_ipo_n80), .B1 (n_0_0_743), .B2 (hfn_ipo_n62));
AOI21_X1 i_0_0_878 (.ZN (n_0_0_756), .A (n_0_0_755), .B1 (n_0_0_717), .B2 (hfn_ipo_n77));
AOI21_X1 i_0_0_877 (.ZN (n_0_0_755), .A (n_0_0_754), .B1 (n_0_0_400), .B2 (drc_ipo_n84));
INV_X1 i_0_0_876 (.ZN (n_0_0_754), .A (n_0_0_733));
NAND2_X1 i_0_0_875 (.ZN (\partialProd[60] ), .A1 (n_0_0_749), .A2 (n_0_0_753));
AOI22_X1 i_0_0_874 (.ZN (n_0_0_753), .A1 (hfn_ipo_n67), .A2 (n_0_0_752), .B1 (hfn_ipo_n71), .B2 (n_0_0_740));
AOI22_X1 i_0_0_873 (.ZN (n_0_0_752), .A1 (n_0_0_751), .A2 (hfn_ipo_n62), .B1 (hfn_ipo_n80), .B2 (n_0_0_729));
AOI21_X1 i_0_0_872 (.ZN (n_0_0_751), .A (n_0_0_750), .B1 (hfn_ipo_n77), .B2 (n_0_0_707));
AOI211_X1 i_0_0_871 (.ZN (n_0_0_750), .A (hfn_ipo_n78), .B (n_0_0_460), .C1 (n_0_0_384), .C2 (drc_ipo_n84));
AOI22_X1 i_0_0_870 (.ZN (n_0_0_749), .A1 (hfn_ipo_n65), .A2 (n_0_0_748), .B1 (hfn_ipo_n69), .B2 (n_0_0_744));
AOI21_X1 i_0_0_869 (.ZN (n_0_0_748), .A (n_0_0_747), .B1 (hfn_ipo_n80), .B2 (n_0_0_734));
AOI221_X1 i_0_0_868 (.ZN (n_0_0_747), .A (hfn_ipo_n80), .B1 (n_0_0_713), .B2 (hfn_ipo_n77)
    , .C1 (n_0_0_746), .C2 (n_0_0_733));
NAND2_X1 i_0_0_867 (.ZN (n_0_0_746), .A1 (n_0_0_393), .A2 (drc_ipo_n84));
NAND2_X1 i_0_0_866 (.ZN (\partialProd[59] ), .A1 (n_0_0_741), .A2 (n_0_0_745));
AOI22_X1 i_0_0_865 (.ZN (n_0_0_745), .A1 (hfn_ipo_n65), .A2 (n_0_0_744), .B1 (hfn_ipo_n69), .B2 (n_0_0_735));
OAI22_X1 i_0_0_864 (.ZN (n_0_0_744), .A1 (n_0_0_718), .A2 (hfn_ipo_n62), .B1 (n_0_0_743), .B2 (hfn_ipo_n80));
AOI22_X1 i_0_0_863 (.ZN (n_0_0_743), .A1 (n_0_0_742), .A2 (n_0_0_733), .B1 (n_0_0_703), .B2 (hfn_ipo_n77));
NAND2_X1 i_0_0_862 (.ZN (n_0_0_742), .A1 (n_0_0_370), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_861 (.ZN (n_0_0_741), .A1 (hfn_ipo_n67), .A2 (n_0_0_740), .B1 (hfn_ipo_n71), .B2 (n_0_0_730));
AOI22_X1 i_0_0_860 (.ZN (n_0_0_740), .A1 (n_0_0_739), .A2 (hfn_ipo_n62), .B1 (n_0_0_724), .B2 (hfn_ipo_n80));
AOI22_X1 i_0_0_859 (.ZN (n_0_0_739), .A1 (n_0_0_738), .A2 (hfn_ipo_n59), .B1 (n_0_0_697), .B2 (hfn_ipo_n77));
INV_X1 i_0_0_858 (.ZN (n_0_0_738), .A (n_0_0_737));
AOI21_X1 i_0_0_857 (.ZN (n_0_0_737), .A (n_0_0_614), .B1 (n_0_0_377), .B2 (drc_ipo_n84));
NAND2_X1 i_0_0_856 (.ZN (\partialProd[58] ), .A1 (n_0_0_731), .A2 (n_0_0_736));
AOI22_X1 i_0_0_855 (.ZN (n_0_0_736), .A1 (hfn_ipo_n65), .A2 (n_0_0_735), .B1 (hfn_ipo_n69), .B2 (n_0_0_719));
OAI22_X1 i_0_0_854 (.ZN (n_0_0_735), .A1 (n_0_0_714), .A2 (hfn_ipo_n62), .B1 (hfn_ipo_n80), .B2 (n_0_0_734));
AOI22_X1 i_0_0_853 (.ZN (n_0_0_734), .A1 (n_0_0_690), .A2 (hfn_ipo_n77), .B1 (n_0_0_732), .B2 (n_0_0_733));
NOR2_X1 i_0_0_852 (.ZN (n_0_0_733), .A1 (n_0_0_631), .A2 (hfn_ipo_n77));
NAND2_X1 i_0_0_851 (.ZN (n_0_0_732), .A1 (n_0_0_353), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_850 (.ZN (n_0_0_731), .A1 (hfn_ipo_n67), .A2 (n_0_0_730), .B1 (hfn_ipo_n71), .B2 (n_0_0_725));
AOI22_X1 i_0_0_849 (.ZN (n_0_0_730), .A1 (n_0_0_708), .A2 (hfn_ipo_n80), .B1 (hfn_ipo_n62), .B2 (n_0_0_729));
AOI22_X1 i_0_0_848 (.ZN (n_0_0_729), .A1 (n_0_0_728), .A2 (hfn_ipo_n59), .B1 (n_0_0_685), .B2 (hfn_ipo_n77));
AOI21_X1 i_0_0_847 (.ZN (n_0_0_728), .A (n_0_0_460), .B1 (n_0_0_727), .B2 (drc_ipo_n84));
INV_X1 i_0_0_846 (.ZN (n_0_0_727), .A (n_0_0_363));
NAND2_X1 i_0_0_845 (.ZN (\partialProd[57] ), .A1 (n_0_0_720), .A2 (n_0_0_726));
AOI22_X1 i_0_0_844 (.ZN (n_0_0_726), .A1 (hfn_ipo_n67), .A2 (n_0_0_725), .B1 (hfn_ipo_n71), .B2 (n_0_0_709));
AOI22_X1 i_0_0_843 (.ZN (n_0_0_725), .A1 (hfn_ipo_n62), .A2 (n_0_0_724), .B1 (n_0_0_698), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_842 (.ZN (n_0_0_724), .A1 (n_0_0_680), .A2 (hfn_ipo_n59), .B1 (n_0_0_723), .B2 (hfn_ipo_n78));
INV_X1 i_0_0_841 (.ZN (n_0_0_723), .A (n_0_0_722));
AOI22_X1 i_0_0_840 (.ZN (n_0_0_722), .A1 (n_0_0_638), .A2 (hfn_ipo_n76), .B1 (n_0_0_721), .B2 (n_0_0_620));
NAND2_X1 i_0_0_839 (.ZN (n_0_0_721), .A1 (n_0_0_345), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_838 (.ZN (n_0_0_720), .A1 (hfn_ipo_n65), .A2 (n_0_0_719), .B1 (hfn_ipo_n69), .B2 (n_0_0_715));
AOI22_X1 i_0_0_837 (.ZN (n_0_0_719), .A1 (n_0_0_704), .A2 (hfn_ipo_n80), .B1 (n_0_0_718), .B2 (hfn_ipo_n62));
AOI22_X1 i_0_0_836 (.ZN (n_0_0_718), .A1 (n_0_0_675), .A2 (hfn_ipo_n77), .B1 (hfn_ipo_n59), .B2 (n_0_0_717));
OAI21_X1 i_0_0_835 (.ZN (n_0_0_717), .A (n_0_0_434), .B1 (n_0_0_338), .B2 (n_0_0_7));
NAND2_X1 i_0_0_834 (.ZN (\partialProd[56] ), .A1 (n_0_0_710), .A2 (n_0_0_716));
AOI22_X1 i_0_0_833 (.ZN (n_0_0_716), .A1 (hfn_ipo_n65), .A2 (n_0_0_715), .B1 (hfn_ipo_n71), .B2 (n_0_0_699));
AOI22_X1 i_0_0_832 (.ZN (n_0_0_715), .A1 (n_0_0_714), .A2 (hfn_ipo_n62), .B1 (n_0_0_691), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_831 (.ZN (n_0_0_714), .A1 (n_0_0_670), .A2 (hfn_ipo_n59), .B1 (hfn_ipo_n77), .B2 (n_0_0_713));
OAI21_X1 i_0_0_830 (.ZN (n_0_0_713), .A (n_0_0_712), .B1 (n_0_0_626), .B2 (hfn_ipo_n73));
OAI21_X1 i_0_0_829 (.ZN (n_0_0_712), .A (n_0_0_632), .B1 (n_0_0_711), .B2 (n_0_0_7));
INV_X1 i_0_0_828 (.ZN (n_0_0_711), .A (n_0_0_322));
AOI22_X1 i_0_0_827 (.ZN (n_0_0_710), .A1 (hfn_ipo_n67), .A2 (n_0_0_709), .B1 (hfn_ipo_n69), .B2 (n_0_0_705));
AOI22_X1 i_0_0_826 (.ZN (n_0_0_709), .A1 (n_0_0_708), .A2 (hfn_ipo_n62), .B1 (hfn_ipo_n80), .B2 (n_0_0_686));
AOI22_X1 i_0_0_825 (.ZN (n_0_0_708), .A1 (n_0_0_665), .A2 (hfn_ipo_n77), .B1 (n_0_0_707), .B2 (hfn_ipo_n59));
OAI21_X1 i_0_0_824 (.ZN (n_0_0_707), .A (n_0_0_425), .B1 (n_0_0_329), .B2 (n_0_0_7));
NAND2_X1 i_0_0_823 (.ZN (\partialProd[55] ), .A1 (n_0_0_700), .A2 (n_0_0_706));
AOI22_X1 i_0_0_822 (.ZN (n_0_0_706), .A1 (hfn_ipo_n65), .A2 (n_0_0_705), .B1 (hfn_ipo_n71), .B2 (n_0_0_687));
AOI22_X1 i_0_0_821 (.ZN (n_0_0_705), .A1 (n_0_0_676), .A2 (hfn_ipo_n80), .B1 (n_0_0_704), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_820 (.ZN (n_0_0_704), .A1 (n_0_0_660), .A2 (hfn_ipo_n59), .B1 (hfn_ipo_n77), .B2 (n_0_0_703));
OAI21_X1 i_0_0_819 (.ZN (n_0_0_703), .A (n_0_0_702), .B1 (hfn_ipo_n73), .B2 (n_0_0_609));
OAI21_X1 i_0_0_818 (.ZN (n_0_0_702), .A (n_0_0_632), .B1 (n_0_0_701), .B2 (n_0_0_7));
INV_X1 i_0_0_817 (.ZN (n_0_0_701), .A (n_0_0_311));
AOI22_X1 i_0_0_816 (.ZN (n_0_0_700), .A1 (hfn_ipo_n67), .A2 (n_0_0_699), .B1 (hfn_ipo_n69), .B2 (n_0_0_692));
AOI22_X1 i_0_0_815 (.ZN (n_0_0_699), .A1 (n_0_0_681), .A2 (hfn_ipo_n80), .B1 (n_0_0_698), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_814 (.ZN (n_0_0_698), .A1 (n_0_0_655), .A2 (hfn_ipo_n59), .B1 (n_0_0_697), .B2 (hfn_ipo_n77));
OAI22_X1 i_0_0_813 (.ZN (n_0_0_697), .A1 (n_0_0_695), .A2 (n_0_0_696), .B1 (n_0_0_615), .B2 (n_0_0_318));
INV_X1 i_0_0_812 (.ZN (n_0_0_696), .A (n_0_0_620));
INV_X1 i_0_0_811 (.ZN (n_0_0_695), .A (n_0_0_694));
NAND2_X1 i_0_0_810 (.ZN (n_0_0_694), .A1 (n_0_0_316), .A2 (drc_ipo_n84));
NAND2_X1 i_0_0_809 (.ZN (\partialProd[54] ), .A1 (n_0_0_688), .A2 (n_0_0_693));
AOI22_X1 i_0_0_808 (.ZN (n_0_0_693), .A1 (hfn_ipo_n65), .A2 (n_0_0_692), .B1 (hfn_ipo_n71), .B2 (n_0_0_682));
AOI22_X1 i_0_0_807 (.ZN (n_0_0_692), .A1 (n_0_0_671), .A2 (hfn_ipo_n80), .B1 (n_0_0_691), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_806 (.ZN (n_0_0_691), .A1 (n_0_0_650), .A2 (hfn_ipo_n59), .B1 (hfn_ipo_n77), .B2 (n_0_0_690));
OAI21_X1 i_0_0_805 (.ZN (n_0_0_690), .A (n_0_0_689), .B1 (n_0_0_604), .B2 (hfn_ipo_n73));
OAI21_X1 i_0_0_804 (.ZN (n_0_0_689), .A (n_0_0_632), .B1 (n_0_0_299), .B2 (n_0_0_7));
AOI22_X1 i_0_0_803 (.ZN (n_0_0_688), .A1 (hfn_ipo_n67), .A2 (n_0_0_687), .B1 (hfn_ipo_n69), .B2 (n_0_0_677));
AOI22_X1 i_0_0_802 (.ZN (n_0_0_687), .A1 (n_0_0_666), .A2 (hfn_ipo_n80), .B1 (hfn_ipo_n62), .B2 (n_0_0_686));
OAI22_X1 i_0_0_801 (.ZN (n_0_0_686), .A1 (n_0_0_645), .A2 (hfn_ipo_n59), .B1 (n_0_0_685), .B2 (hfn_ipo_n77));
OAI21_X1 i_0_0_800 (.ZN (n_0_0_685), .A (n_0_0_684), .B1 (n_0_0_597), .B2 (hfn_ipo_n73));
OAI21_X1 i_0_0_799 (.ZN (n_0_0_684), .A (n_0_0_620), .B1 (n_0_0_306), .B2 (n_0_0_7));
NAND2_X1 i_0_0_798 (.ZN (\partialProd[53] ), .A1 (n_0_0_678), .A2 (n_0_0_683));
AOI22_X1 i_0_0_797 (.ZN (n_0_0_683), .A1 (hfn_ipo_n67), .A2 (n_0_0_682), .B1 (hfn_ipo_n71), .B2 (n_0_0_667));
AOI22_X1 i_0_0_796 (.ZN (n_0_0_682), .A1 (n_0_0_656), .A2 (hfn_ipo_n80), .B1 (hfn_ipo_n62), .B2 (n_0_0_681));
OAI22_X1 i_0_0_795 (.ZN (n_0_0_681), .A1 (n_0_0_640), .A2 (hfn_ipo_n59), .B1 (n_0_0_680), .B2 (hfn_ipo_n78));
OAI21_X1 i_0_0_794 (.ZN (n_0_0_680), .A (n_0_0_679), .B1 (n_0_0_591), .B2 (n_0_0_318));
OAI21_X1 i_0_0_793 (.ZN (n_0_0_679), .A (n_0_0_620), .B1 (n_0_0_284), .B2 (n_0_0_7));
AOI22_X1 i_0_0_792 (.ZN (n_0_0_678), .A1 (hfn_ipo_n65), .A2 (n_0_0_677), .B1 (hfn_ipo_n69), .B2 (n_0_0_672));
AOI22_X1 i_0_0_791 (.ZN (n_0_0_677), .A1 (n_0_0_661), .A2 (hfn_ipo_n80), .B1 (n_0_0_676), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_790 (.ZN (n_0_0_676), .A1 (n_0_0_634), .A2 (hfn_ipo_n59), .B1 (n_0_0_675), .B2 (hfn_ipo_n77));
OAI21_X1 i_0_0_789 (.ZN (n_0_0_675), .A (n_0_0_674), .B1 (n_0_0_585), .B2 (hfn_ipo_n73));
OAI21_X1 i_0_0_788 (.ZN (n_0_0_674), .A (n_0_0_632), .B1 (n_0_0_292), .B2 (n_0_0_7));
NAND2_X1 i_0_0_787 (.ZN (\partialProd[52] ), .A1 (n_0_0_668), .A2 (n_0_0_673));
AOI22_X1 i_0_0_786 (.ZN (n_0_0_673), .A1 (hfn_ipo_n65), .A2 (n_0_0_672), .B1 (hfn_ipo_n71), .B2 (n_0_0_657));
AOI22_X1 i_0_0_785 (.ZN (n_0_0_672), .A1 (n_0_0_651), .A2 (hfn_ipo_n80), .B1 (n_0_0_671), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_784 (.ZN (n_0_0_671), .A1 (n_0_0_627), .A2 (hfn_ipo_n59), .B1 (n_0_0_670), .B2 (hfn_ipo_n77));
OAI21_X1 i_0_0_783 (.ZN (n_0_0_670), .A (n_0_0_669), .B1 (n_0_0_580), .B2 (hfn_ipo_n73));
OAI21_X1 i_0_0_782 (.ZN (n_0_0_669), .A (n_0_0_632), .B1 (n_0_0_390), .B2 (n_0_0_7));
AOI22_X1 i_0_0_781 (.ZN (n_0_0_668), .A1 (hfn_ipo_n67), .A2 (n_0_0_667), .B1 (hfn_ipo_n69), .B2 (n_0_0_662));
AOI22_X1 i_0_0_780 (.ZN (n_0_0_667), .A1 (n_0_0_666), .A2 (hfn_ipo_n62), .B1 (n_0_0_646), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_779 (.ZN (n_0_0_666), .A1 (n_0_0_665), .A2 (hfn_ipo_n77), .B1 (n_0_0_622), .B2 (hfn_ipo_n59));
AOI222_X1 i_0_0_778 (.ZN (n_0_0_665), .A1 (n_0_0_575), .A2 (hfn_ipo_n75), .B1 (n_0_0_47)
    , .B2 (n_0_0_277), .C1 (n_0_0_664), .C2 (n_0_0_10));
INV_X1 i_0_0_777 (.ZN (n_0_0_664), .A (\extended_M[63] ));
NAND2_X1 i_0_0_776 (.ZN (\partialProd[51] ), .A1 (n_0_0_658), .A2 (n_0_0_663));
AOI22_X1 i_0_0_775 (.ZN (n_0_0_663), .A1 (hfn_ipo_n65), .A2 (n_0_0_662), .B1 (hfn_ipo_n69), .B2 (n_0_0_652));
AOI22_X1 i_0_0_774 (.ZN (n_0_0_662), .A1 (n_0_0_635), .A2 (hfn_ipo_n80), .B1 (n_0_0_661), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_773 (.ZN (n_0_0_661), .A1 (n_0_0_610), .A2 (hfn_ipo_n59), .B1 (n_0_0_660), .B2 (hfn_ipo_n77));
OAI21_X1 i_0_0_772 (.ZN (n_0_0_660), .A (n_0_0_659), .B1 (n_0_0_563), .B2 (hfn_ipo_n73));
OAI21_X1 i_0_0_771 (.ZN (n_0_0_659), .A (n_0_0_632), .B1 (n_0_0_367), .B2 (n_0_0_7));
AOI22_X1 i_0_0_770 (.ZN (n_0_0_658), .A1 (hfn_ipo_n67), .A2 (n_0_0_657), .B1 (hfn_ipo_n71), .B2 (n_0_0_647));
AOI22_X1 i_0_0_769 (.ZN (n_0_0_657), .A1 (n_0_0_641), .A2 (hfn_ipo_n80), .B1 (n_0_0_656), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_768 (.ZN (n_0_0_656), .A1 (n_0_0_616), .A2 (hfn_ipo_n59), .B1 (n_0_0_655), .B2 (hfn_ipo_n78));
OAI21_X1 i_0_0_767 (.ZN (n_0_0_655), .A (n_0_0_654), .B1 (n_0_0_569), .B2 (n_0_0_318));
OAI21_X1 i_0_0_766 (.ZN (n_0_0_654), .A (n_0_0_620), .B1 (n_0_0_265), .B2 (n_0_0_7));
NAND2_X1 i_0_0_765 (.ZN (\partialProd[50] ), .A1 (n_0_0_648), .A2 (n_0_0_653));
AOI22_X1 i_0_0_764 (.ZN (n_0_0_653), .A1 (hfn_ipo_n65), .A2 (n_0_0_652), .B1 (hfn_ipo_n69), .B2 (n_0_0_636));
OAI22_X1 i_0_0_763 (.ZN (n_0_0_652), .A1 (n_0_0_628), .A2 (hfn_ipo_n62), .B1 (n_0_0_651), .B2 (hfn_ipo_n80));
AOI22_X1 i_0_0_762 (.ZN (n_0_0_651), .A1 (n_0_0_605), .A2 (hfn_ipo_n77), .B1 (n_0_0_650), .B2 (hfn_ipo_n59));
OAI21_X1 i_0_0_761 (.ZN (n_0_0_650), .A (n_0_0_649), .B1 (n_0_0_558), .B2 (hfn_ipo_n73));
OAI21_X1 i_0_0_760 (.ZN (n_0_0_649), .A (n_0_0_632), .B1 (n_0_0_350), .B2 (n_0_0_603));
AOI22_X1 i_0_0_759 (.ZN (n_0_0_648), .A1 (hfn_ipo_n67), .A2 (n_0_0_647), .B1 (hfn_ipo_n71), .B2 (n_0_0_642));
AOI22_X1 i_0_0_758 (.ZN (n_0_0_647), .A1 (n_0_0_646), .A2 (hfn_ipo_n62), .B1 (n_0_0_623), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_757 (.ZN (n_0_0_646), .A1 (n_0_0_598), .A2 (hfn_ipo_n59), .B1 (hfn_ipo_n77), .B2 (n_0_0_645));
OAI21_X1 i_0_0_756 (.ZN (n_0_0_645), .A (n_0_0_644), .B1 (n_0_0_553), .B2 (n_0_0_318));
OAI21_X1 i_0_0_755 (.ZN (n_0_0_644), .A (n_0_0_620), .B1 (n_0_0_248), .B2 (n_0_0_7));
NAND2_X1 i_0_0_754 (.ZN (\partialProd[49] ), .A1 (n_0_0_637), .A2 (n_0_0_643));
AOI22_X1 i_0_0_753 (.ZN (n_0_0_643), .A1 (hfn_ipo_n67), .A2 (n_0_0_642), .B1 (hfn_ipo_n71), .B2 (n_0_0_624));
OAI22_X1 i_0_0_752 (.ZN (n_0_0_642), .A1 (n_0_0_641), .A2 (hfn_ipo_n80), .B1 (n_0_0_617), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_751 (.ZN (n_0_0_641), .A1 (n_0_0_592), .A2 (hfn_ipo_n59), .B1 (hfn_ipo_n78), .B2 (n_0_0_640));
OAI22_X1 i_0_0_750 (.ZN (n_0_0_640), .A1 (n_0_0_639), .A2 (hfn_ipo_n76), .B1 (n_0_0_547), .B2 (n_0_0_318));
INV_X1 i_0_0_749 (.ZN (n_0_0_639), .A (n_0_0_638));
AOI21_X1 i_0_0_748 (.ZN (n_0_0_638), .A (n_0_0_460), .B1 (n_0_0_240), .B2 (drc_ipo_n84));
AOI22_X1 i_0_0_747 (.ZN (n_0_0_637), .A1 (hfn_ipo_n65), .A2 (n_0_0_636), .B1 (hfn_ipo_n69), .B2 (n_0_0_629));
AOI22_X1 i_0_0_746 (.ZN (n_0_0_636), .A1 (n_0_0_611), .A2 (hfn_ipo_n80), .B1 (n_0_0_635), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_745 (.ZN (n_0_0_635), .A1 (n_0_0_586), .A2 (hfn_ipo_n59), .B1 (n_0_0_634), .B2 (hfn_ipo_n77));
OAI21_X1 i_0_0_744 (.ZN (n_0_0_634), .A (n_0_0_633), .B1 (n_0_0_541), .B2 (hfn_ipo_n73));
OAI21_X1 i_0_0_743 (.ZN (n_0_0_633), .A (n_0_0_632), .B1 (n_0_0_234), .B2 (n_0_0_7));
NOR2_X1 i_0_0_742 (.ZN (n_0_0_632), .A1 (n_0_0_631), .A2 (hfn_ipo_n75));
NOR2_X1 i_0_0_741 (.ZN (n_0_0_631), .A1 (\extended_M_mul_neg_one[63] ), .A2 (drc_ipo_n84));
NAND2_X1 i_0_0_740 (.ZN (\partialProd[48] ), .A1 (n_0_0_625), .A2 (n_0_0_630));
AOI22_X1 i_0_0_739 (.ZN (n_0_0_630), .A1 (hfn_ipo_n65), .A2 (n_0_0_629), .B1 (hfn_ipo_n69), .B2 (n_0_0_612));
OAI22_X1 i_0_0_738 (.ZN (n_0_0_629), .A1 (n_0_0_606), .A2 (hfn_ipo_n62), .B1 (n_0_0_628), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_737 (.ZN (n_0_0_628), .A1 (n_0_0_581), .A2 (hfn_ipo_n59), .B1 (n_0_0_627), .B2 (hfn_ipo_n77));
OAI22_X1 i_0_0_736 (.ZN (n_0_0_627), .A1 (n_0_0_536), .A2 (hfn_ipo_n73), .B1 (hfn_ipo_n75), .B2 (n_0_0_626));
AOI21_X1 i_0_0_735 (.ZN (n_0_0_626), .A (n_0_0_603), .B1 (n_0_0_227), .B2 (drc_ipo_n84));
AOI22_X1 i_0_0_734 (.ZN (n_0_0_625), .A1 (hfn_ipo_n67), .A2 (n_0_0_624), .B1 (hfn_ipo_n71), .B2 (n_0_0_618));
AOI22_X1 i_0_0_733 (.ZN (n_0_0_624), .A1 (n_0_0_599), .A2 (hfn_ipo_n80), .B1 (n_0_0_623), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_732 (.ZN (n_0_0_623), .A1 (n_0_0_576), .A2 (hfn_ipo_n59), .B1 (hfn_ipo_n77), .B2 (n_0_0_622));
OAI21_X1 i_0_0_731 (.ZN (n_0_0_622), .A (n_0_0_621), .B1 (n_0_0_531), .B2 (n_0_0_318));
OAI21_X1 i_0_0_730 (.ZN (n_0_0_621), .A (n_0_0_620), .B1 (n_0_0_220), .B2 (n_0_0_7));
NOR2_X1 i_0_0_729 (.ZN (n_0_0_620), .A1 (n_0_0_460), .A2 (hfn_ipo_n76));
NAND2_X1 i_0_0_728 (.ZN (\partialProd[47] ), .A1 (n_0_0_613), .A2 (n_0_0_619));
AOI22_X1 i_0_0_727 (.ZN (n_0_0_619), .A1 (hfn_ipo_n67), .A2 (n_0_0_618), .B1 (hfn_ipo_n69), .B2 (n_0_0_607));
AOI22_X1 i_0_0_726 (.ZN (n_0_0_618), .A1 (n_0_0_593), .A2 (hfn_ipo_n80), .B1 (n_0_0_617), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_725 (.ZN (n_0_0_617), .A1 (n_0_0_616), .A2 (hfn_ipo_n78), .B1 (n_0_0_570), .B2 (hfn_ipo_n60));
AOI22_X1 i_0_0_724 (.ZN (n_0_0_616), .A1 (n_0_0_520), .A2 (hfn_ipo_n76), .B1 (n_0_0_318), .B2 (n_0_0_615));
AOI21_X1 i_0_0_723 (.ZN (n_0_0_615), .A (n_0_0_614), .B1 (n_0_0_442), .B2 (\extended_M[15] ));
INV_X1 i_0_0_722 (.ZN (n_0_0_614), .A (n_0_0_425));
AOI22_X1 i_0_0_721 (.ZN (n_0_0_613), .A1 (hfn_ipo_n65), .A2 (n_0_0_612), .B1 (hfn_ipo_n71), .B2 (n_0_0_600));
AOI22_X1 i_0_0_720 (.ZN (n_0_0_612), .A1 (n_0_0_587), .A2 (hfn_ipo_n80), .B1 (n_0_0_611), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_719 (.ZN (n_0_0_611), .A1 (n_0_0_564), .A2 (hfn_ipo_n59), .B1 (n_0_0_610), .B2 (hfn_ipo_n77));
AOI22_X1 i_0_0_718 (.ZN (n_0_0_610), .A1 (n_0_0_525), .A2 (hfn_ipo_n75), .B1 (hfn_ipo_n73), .B2 (n_0_0_609));
AOI21_X1 i_0_0_717 (.ZN (n_0_0_609), .A (n_0_0_603), .B1 (n_0_0_442), .B2 (\extended_M_mul_neg_one[15] ));
NAND2_X1 i_0_0_716 (.ZN (\partialProd[46] ), .A1 (n_0_0_601), .A2 (n_0_0_608));
AOI22_X1 i_0_0_715 (.ZN (n_0_0_608), .A1 (hfn_ipo_n65), .A2 (n_0_0_607), .B1 (hfn_ipo_n71), .B2 (n_0_0_594));
OAI22_X1 i_0_0_714 (.ZN (n_0_0_607), .A1 (n_0_0_582), .A2 (hfn_ipo_n62), .B1 (n_0_0_606), .B2 (hfn_ipo_n80));
AOI22_X1 i_0_0_713 (.ZN (n_0_0_606), .A1 (n_0_0_559), .A2 (hfn_ipo_n77), .B1 (n_0_0_605), .B2 (hfn_ipo_n59));
OAI22_X1 i_0_0_712 (.ZN (n_0_0_605), .A1 (n_0_0_515), .A2 (hfn_ipo_n73), .B1 (n_0_0_604), .B2 (hfn_ipo_n75));
OAI22_X1 i_0_0_711 (.ZN (n_0_0_604), .A1 (n_0_0_602), .A2 (n_0_0_603), .B1 (n_0_0_411), .B2 (n_0_0_15));
INV_X1 i_0_0_710 (.ZN (n_0_0_603), .A (n_0_0_434));
OAI21_X1 i_0_0_709 (.ZN (n_0_0_602), .A (n_0_0_15), .B1 (n_0_0_197), .B2 (n_0_0_7));
AOI22_X1 i_0_0_708 (.ZN (n_0_0_601), .A1 (hfn_ipo_n67), .A2 (n_0_0_600), .B1 (hfn_ipo_n69), .B2 (n_0_0_588));
AOI22_X1 i_0_0_707 (.ZN (n_0_0_600), .A1 (n_0_0_577), .A2 (hfn_ipo_n80), .B1 (n_0_0_599), .B2 (hfn_ipo_n62));
OAI22_X1 i_0_0_706 (.ZN (n_0_0_599), .A1 (n_0_0_598), .A2 (hfn_ipo_n77), .B1 (hfn_ipo_n59), .B2 (n_0_0_554));
OAI22_X1 i_0_0_705 (.ZN (n_0_0_598), .A1 (n_0_0_510), .A2 (hfn_ipo_n73), .B1 (hfn_ipo_n75), .B2 (n_0_0_597));
AOI22_X1 i_0_0_704 (.ZN (n_0_0_597), .A1 (n_0_0_461), .A2 (n_0_0_596), .B1 (\extended_M[30] ), .B2 (n_0_0_412));
OR2_X1 i_0_0_703 (.ZN (n_0_0_596), .A1 (n_0_0_7), .A2 (\extended_M[14] ));
NAND2_X1 i_0_0_702 (.ZN (\partialProd[45] ), .A1 (n_0_0_589), .A2 (n_0_0_595));
AOI22_X1 i_0_0_701 (.ZN (n_0_0_595), .A1 (hfn_ipo_n67), .A2 (n_0_0_594), .B1 (hfn_ipo_n71), .B2 (n_0_0_578));
AOI22_X1 i_0_0_700 (.ZN (n_0_0_594), .A1 (n_0_0_593), .A2 (hfn_ipo_n63), .B1 (n_0_0_571), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_699 (.ZN (n_0_0_593), .A1 (n_0_0_592), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_548));
AOI22_X1 i_0_0_698 (.ZN (n_0_0_592), .A1 (n_0_0_505), .A2 (hfn_ipo_n76), .B1 (n_0_0_318), .B2 (n_0_0_591));
AOI22_X1 i_0_0_697 (.ZN (n_0_0_591), .A1 (n_0_0_461), .A2 (n_0_0_590), .B1 (\extended_M[29] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_696 (.ZN (n_0_0_590), .A1 (n_0_0_186), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_695 (.ZN (n_0_0_589), .A1 (hfn_ipo_n65), .A2 (n_0_0_588), .B1 (hfn_ipo_n69), .B2 (n_0_0_583));
AOI22_X1 i_0_0_694 (.ZN (n_0_0_588), .A1 (n_0_0_587), .A2 (hfn_ipo_n62), .B1 (n_0_0_565), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_693 (.ZN (n_0_0_587), .A1 (n_0_0_586), .A2 (hfn_ipo_n77), .B1 (n_0_0_542), .B2 (hfn_ipo_n59));
AOI22_X1 i_0_0_692 (.ZN (n_0_0_586), .A1 (n_0_0_500), .A2 (hfn_ipo_n75), .B1 (n_0_0_585), .B2 (hfn_ipo_n73));
AOI221_X1 i_0_0_691 (.ZN (n_0_0_585), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[13] )
    , .B2 (n_0_0_442), .C1 (\extended_M_mul_neg_one[29] ), .C2 (n_0_0_412));
NAND2_X1 i_0_0_690 (.ZN (\partialProd[44] ), .A1 (n_0_0_579), .A2 (n_0_0_584));
AOI22_X1 i_0_0_689 (.ZN (n_0_0_584), .A1 (hfn_ipo_n65), .A2 (n_0_0_583), .B1 (hfn_ipo_n69), .B2 (n_0_0_566));
AOI22_X1 i_0_0_688 (.ZN (n_0_0_583), .A1 (n_0_0_582), .A2 (hfn_ipo_n62), .B1 (n_0_0_560), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_687 (.ZN (n_0_0_582), .A1 (n_0_0_581), .A2 (hfn_ipo_n77), .B1 (n_0_0_537), .B2 (hfn_ipo_n59));
OAI22_X1 i_0_0_686 (.ZN (n_0_0_581), .A1 (n_0_0_490), .A2 (hfn_ipo_n73), .B1 (n_0_0_580), .B2 (hfn_ipo_n75));
AOI221_X1 i_0_0_685 (.ZN (n_0_0_580), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[28] )
    , .B2 (n_0_0_412), .C1 (\extended_M_mul_neg_one[12] ), .C2 (n_0_0_442));
AOI22_X1 i_0_0_684 (.ZN (n_0_0_579), .A1 (hfn_ipo_n67), .A2 (n_0_0_578), .B1 (hfn_ipo_n71), .B2 (n_0_0_572));
AOI22_X1 i_0_0_683 (.ZN (n_0_0_578), .A1 (n_0_0_577), .A2 (hfn_ipo_n62), .B1 (n_0_0_555), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_682 (.ZN (n_0_0_577), .A1 (n_0_0_576), .A2 (hfn_ipo_n77), .B1 (n_0_0_532), .B2 (hfn_ipo_n59));
AOI22_X1 i_0_0_681 (.ZN (n_0_0_576), .A1 (n_0_0_495), .A2 (hfn_ipo_n75), .B1 (n_0_0_575), .B2 (hfn_ipo_n73));
AOI22_X1 i_0_0_680 (.ZN (n_0_0_575), .A1 (n_0_0_461), .A2 (n_0_0_574), .B1 (\extended_M[28] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_679 (.ZN (n_0_0_574), .A1 (n_0_0_180), .A2 (drc_ipo_n84));
NAND2_X1 i_0_0_678 (.ZN (\partialProd[43] ), .A1 (n_0_0_567), .A2 (n_0_0_573));
AOI22_X1 i_0_0_677 (.ZN (n_0_0_573), .A1 (hfn_ipo_n67), .A2 (n_0_0_572), .B1 (hfn_ipo_n69), .B2 (n_0_0_561));
AOI22_X1 i_0_0_676 (.ZN (n_0_0_572), .A1 (n_0_0_549), .A2 (hfn_ipo_n81), .B1 (n_0_0_571), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_675 (.ZN (n_0_0_571), .A1 (n_0_0_521), .A2 (hfn_ipo_n60), .B1 (hfn_ipo_n78), .B2 (n_0_0_570));
AOI22_X1 i_0_0_674 (.ZN (n_0_0_570), .A1 (n_0_0_480), .A2 (hfn_ipo_n76), .B1 (n_0_0_569), .B2 (n_0_0_318));
AOI22_X1 i_0_0_673 (.ZN (n_0_0_569), .A1 (n_0_0_461), .A2 (n_0_0_568), .B1 (\extended_M[27] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_672 (.ZN (n_0_0_568), .A1 (n_0_0_163), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_671 (.ZN (n_0_0_567), .A1 (hfn_ipo_n65), .A2 (n_0_0_566), .B1 (hfn_ipo_n71), .B2 (n_0_0_556));
AOI22_X1 i_0_0_670 (.ZN (n_0_0_566), .A1 (hfn_ipo_n62), .A2 (n_0_0_565), .B1 (n_0_0_543), .B2 (hfn_ipo_n80));
OAI22_X1 i_0_0_669 (.ZN (n_0_0_565), .A1 (n_0_0_564), .A2 (hfn_ipo_n77), .B1 (n_0_0_526), .B2 (hfn_ipo_n59));
AOI22_X1 i_0_0_668 (.ZN (n_0_0_564), .A1 (n_0_0_485), .A2 (hfn_ipo_n75), .B1 (n_0_0_563), .B2 (hfn_ipo_n73));
AOI221_X1 i_0_0_667 (.ZN (n_0_0_563), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[27] )
    , .B2 (n_0_0_412), .C1 (\extended_M_mul_neg_one[11] ), .C2 (n_0_0_442));
NAND2_X1 i_0_0_666 (.ZN (\partialProd[42] ), .A1 (n_0_0_557), .A2 (n_0_0_562));
AOI22_X1 i_0_0_665 (.ZN (n_0_0_562), .A1 (hfn_ipo_n65), .A2 (n_0_0_561), .B1 (hfn_ipo_n69), .B2 (n_0_0_544));
AOI22_X1 i_0_0_664 (.ZN (n_0_0_561), .A1 (n_0_0_538), .A2 (hfn_ipo_n81), .B1 (n_0_0_560), .B2 (hfn_ipo_n63));
AOI22_X1 i_0_0_663 (.ZN (n_0_0_560), .A1 (n_0_0_559), .A2 (hfn_ipo_n59), .B1 (n_0_0_516), .B2 (hfn_ipo_n77));
AOI22_X1 i_0_0_662 (.ZN (n_0_0_559), .A1 (n_0_0_558), .A2 (hfn_ipo_n73), .B1 (n_0_0_468), .B2 (hfn_ipo_n75));
AOI221_X1 i_0_0_661 (.ZN (n_0_0_558), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[26] )
    , .B2 (n_0_0_412), .C1 (\extended_M_mul_neg_one[10] ), .C2 (n_0_0_442));
AOI22_X1 i_0_0_660 (.ZN (n_0_0_557), .A1 (hfn_ipo_n67), .A2 (n_0_0_556), .B1 (hfn_ipo_n71), .B2 (n_0_0_550));
AOI22_X1 i_0_0_659 (.ZN (n_0_0_556), .A1 (n_0_0_533), .A2 (hfn_ipo_n81), .B1 (n_0_0_555), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_658 (.ZN (n_0_0_555), .A1 (n_0_0_511), .A2 (hfn_ipo_n59), .B1 (hfn_ipo_n77), .B2 (n_0_0_554));
AOI22_X1 i_0_0_657 (.ZN (n_0_0_554), .A1 (n_0_0_474), .A2 (hfn_ipo_n76), .B1 (n_0_0_553), .B2 (n_0_0_318));
AOI22_X1 i_0_0_656 (.ZN (n_0_0_553), .A1 (n_0_0_461), .A2 (n_0_0_552), .B1 (\extended_M[26] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_655 (.ZN (n_0_0_552), .A1 (n_0_0_153), .A2 (drc_ipo_n84));
NAND2_X1 i_0_0_654 (.ZN (\partialProd[41] ), .A1 (n_0_0_545), .A2 (n_0_0_551));
AOI22_X1 i_0_0_653 (.ZN (n_0_0_551), .A1 (hfn_ipo_n67), .A2 (n_0_0_550), .B1 (hfn_ipo_n69), .B2 (n_0_0_539));
AOI22_X1 i_0_0_652 (.ZN (n_0_0_550), .A1 (n_0_0_549), .A2 (hfn_ipo_n63), .B1 (n_0_0_522), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_651 (.ZN (n_0_0_549), .A1 (n_0_0_506), .A2 (hfn_ipo_n60), .B1 (hfn_ipo_n78), .B2 (n_0_0_548));
AOI22_X1 i_0_0_650 (.ZN (n_0_0_548), .A1 (n_0_0_547), .A2 (n_0_0_318), .B1 (n_0_0_463), .B2 (hfn_ipo_n76));
AOI22_X1 i_0_0_649 (.ZN (n_0_0_547), .A1 (n_0_0_461), .A2 (n_0_0_546), .B1 (\extended_M[25] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_648 (.ZN (n_0_0_546), .A1 (n_0_0_148), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_647 (.ZN (n_0_0_545), .A1 (hfn_ipo_n65), .A2 (n_0_0_544), .B1 (hfn_ipo_n71), .B2 (n_0_0_534));
OAI22_X1 i_0_0_646 (.ZN (n_0_0_544), .A1 (n_0_0_543), .A2 (hfn_ipo_n81), .B1 (n_0_0_527), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_645 (.ZN (n_0_0_543), .A1 (n_0_0_542), .A2 (hfn_ipo_n77), .B1 (n_0_0_501), .B2 (hfn_ipo_n59));
OAI22_X1 i_0_0_644 (.ZN (n_0_0_542), .A1 (n_0_0_455), .A2 (n_0_0_318), .B1 (n_0_0_541), .B2 (hfn_ipo_n75));
AOI221_X1 i_0_0_643 (.ZN (n_0_0_541), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[25] )
    , .B2 (n_0_0_412), .C1 (\extended_M_mul_neg_one[9] ), .C2 (n_0_0_442));
NAND2_X1 i_0_0_642 (.ZN (\partialProd[40] ), .A1 (n_0_0_535), .A2 (n_0_0_540));
AOI22_X1 i_0_0_641 (.ZN (n_0_0_540), .A1 (hfn_ipo_n65), .A2 (n_0_0_539), .B1 (hfn_ipo_n69), .B2 (n_0_0_528));
AOI22_X1 i_0_0_640 (.ZN (n_0_0_539), .A1 (n_0_0_538), .A2 (hfn_ipo_n63), .B1 (n_0_0_517), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_639 (.ZN (n_0_0_538), .A1 (n_0_0_537), .A2 (hfn_ipo_n77), .B1 (n_0_0_491), .B2 (hfn_ipo_n59));
AOI22_X1 i_0_0_638 (.ZN (n_0_0_537), .A1 (n_0_0_536), .A2 (hfn_ipo_n73), .B1 (n_0_0_444), .B2 (hfn_ipo_n75));
AOI221_X1 i_0_0_637 (.ZN (n_0_0_536), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[24] )
    , .B2 (n_0_0_412), .C1 (\extended_M_mul_neg_one[8] ), .C2 (n_0_0_442));
AOI22_X1 i_0_0_636 (.ZN (n_0_0_535), .A1 (hfn_ipo_n67), .A2 (n_0_0_534), .B1 (hfn_ipo_n71), .B2 (n_0_0_523));
AOI22_X1 i_0_0_635 (.ZN (n_0_0_534), .A1 (n_0_0_533), .A2 (hfn_ipo_n63), .B1 (n_0_0_512), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_634 (.ZN (n_0_0_533), .A1 (n_0_0_496), .A2 (hfn_ipo_n60), .B1 (n_0_0_532), .B2 (hfn_ipo_n78));
AOI22_X1 i_0_0_633 (.ZN (n_0_0_532), .A1 (n_0_0_449), .A2 (hfn_ipo_n76), .B1 (n_0_0_318), .B2 (n_0_0_531));
AOI22_X1 i_0_0_632 (.ZN (n_0_0_531), .A1 (n_0_0_461), .A2 (n_0_0_530), .B1 (\extended_M[24] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_631 (.ZN (n_0_0_530), .A1 (n_0_0_135), .A2 (drc_ipo_n84));
NAND2_X1 i_0_0_630 (.ZN (\partialProd[39] ), .A1 (n_0_0_524), .A2 (n_0_0_529));
AOI22_X1 i_0_0_629 (.ZN (n_0_0_529), .A1 (hfn_ipo_n65), .A2 (n_0_0_528), .B1 (hfn_ipo_n71), .B2 (n_0_0_513));
AOI22_X1 i_0_0_628 (.ZN (n_0_0_528), .A1 (n_0_0_502), .A2 (hfn_ipo_n81), .B1 (n_0_0_527), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_627 (.ZN (n_0_0_527), .A1 (n_0_0_486), .A2 (hfn_ipo_n60), .B1 (n_0_0_526), .B2 (hfn_ipo_n78));
AOI22_X1 i_0_0_626 (.ZN (n_0_0_526), .A1 (n_0_0_525), .A2 (n_0_0_318), .B1 (hfn_ipo_n75), .B2 (n_0_0_436));
AOI221_X1 i_0_0_625 (.ZN (n_0_0_525), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[7] )
    , .B2 (n_0_0_442), .C1 (\extended_M_mul_neg_one[23] ), .C2 (n_0_0_412));
AOI22_X1 i_0_0_624 (.ZN (n_0_0_524), .A1 (hfn_ipo_n67), .A2 (n_0_0_523), .B1 (hfn_ipo_n69), .B2 (n_0_0_518));
AOI22_X1 i_0_0_623 (.ZN (n_0_0_523), .A1 (n_0_0_507), .A2 (hfn_ipo_n81), .B1 (n_0_0_522), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_622 (.ZN (n_0_0_522), .A1 (n_0_0_521), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_481));
AOI22_X1 i_0_0_621 (.ZN (n_0_0_521), .A1 (n_0_0_520), .A2 (n_0_0_318), .B1 (hfn_ipo_n76), .B2 (n_0_0_427));
AOI221_X1 i_0_0_620 (.ZN (n_0_0_520), .A (n_0_0_426), .B1 (\extended_M[23] ), .B2 (n_0_0_412)
    , .C1 (\extended_M[7] ), .C2 (n_0_0_442));
NAND2_X1 i_0_0_619 (.ZN (\partialProd[38] ), .A1 (n_0_0_514), .A2 (n_0_0_519));
AOI22_X1 i_0_0_618 (.ZN (n_0_0_519), .A1 (hfn_ipo_n65), .A2 (n_0_0_518), .B1 (hfn_ipo_n71), .B2 (n_0_0_508));
AOI22_X1 i_0_0_617 (.ZN (n_0_0_518), .A1 (hfn_ipo_n63), .A2 (n_0_0_517), .B1 (n_0_0_492), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_616 (.ZN (n_0_0_517), .A1 (n_0_0_469), .A2 (hfn_ipo_n59), .B1 (n_0_0_516), .B2 (hfn_ipo_n78));
AOI22_X1 i_0_0_615 (.ZN (n_0_0_516), .A1 (n_0_0_515), .A2 (hfn_ipo_n73), .B1 (hfn_ipo_n75), .B2 (n_0_0_413));
AOI221_X1 i_0_0_614 (.ZN (n_0_0_515), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[22] )
    , .B2 (n_0_0_412), .C1 (\extended_M_mul_neg_one[6] ), .C2 (n_0_0_442));
AOI22_X1 i_0_0_613 (.ZN (n_0_0_514), .A1 (hfn_ipo_n67), .A2 (n_0_0_513), .B1 (hfn_ipo_n69), .B2 (n_0_0_503));
AOI22_X1 i_0_0_612 (.ZN (n_0_0_513), .A1 (n_0_0_497), .A2 (hfn_ipo_n81), .B1 (n_0_0_512), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_611 (.ZN (n_0_0_512), .A1 (n_0_0_511), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_475));
OAI22_X1 i_0_0_610 (.ZN (n_0_0_511), .A1 (n_0_0_510), .A2 (hfn_ipo_n75), .B1 (n_0_0_8), .B2 (n_0_0_419));
AOI221_X1 i_0_0_609 (.ZN (n_0_0_510), .A (n_0_0_426), .B1 (\extended_M[22] ), .B2 (n_0_0_412)
    , .C1 (\extended_M[6] ), .C2 (n_0_0_442));
NAND2_X1 i_0_0_608 (.ZN (\partialProd[37] ), .A1 (n_0_0_504), .A2 (n_0_0_509));
AOI22_X1 i_0_0_607 (.ZN (n_0_0_509), .A1 (hfn_ipo_n67), .A2 (n_0_0_508), .B1 (hfn_ipo_n69), .B2 (n_0_0_493));
AOI22_X1 i_0_0_606 (.ZN (n_0_0_508), .A1 (n_0_0_507), .A2 (hfn_ipo_n63), .B1 (n_0_0_482), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_605 (.ZN (n_0_0_507), .A1 (n_0_0_506), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_464));
OAI22_X1 i_0_0_604 (.ZN (n_0_0_506), .A1 (n_0_0_505), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_405));
AOI221_X1 i_0_0_603 (.ZN (n_0_0_505), .A (n_0_0_426), .B1 (\extended_M[21] ), .B2 (n_0_0_412)
    , .C1 (\extended_M[5] ), .C2 (n_0_0_442));
AOI22_X1 i_0_0_602 (.ZN (n_0_0_504), .A1 (hfn_ipo_n65), .A2 (n_0_0_503), .B1 (hfn_ipo_n71), .B2 (n_0_0_498));
AOI22_X1 i_0_0_601 (.ZN (n_0_0_503), .A1 (n_0_0_502), .A2 (hfn_ipo_n63), .B1 (n_0_0_487), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_600 (.ZN (n_0_0_502), .A1 (n_0_0_501), .A2 (hfn_ipo_n78), .B1 (n_0_0_456), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_599 (.ZN (n_0_0_501), .A1 (n_0_0_500), .A2 (hfn_ipo_n75), .B1 (n_0_0_8), .B2 (n_0_0_398));
AOI221_X1 i_0_0_598 (.ZN (n_0_0_500), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[21] )
    , .B2 (n_0_0_412), .C1 (\extended_M_mul_neg_one[5] ), .C2 (n_0_0_442));
NAND2_X1 i_0_0_597 (.ZN (\partialProd[36] ), .A1 (n_0_0_494), .A2 (n_0_0_499));
AOI22_X1 i_0_0_596 (.ZN (n_0_0_499), .A1 (hfn_ipo_n67), .A2 (n_0_0_498), .B1 (hfn_ipo_n71), .B2 (n_0_0_483));
AOI22_X1 i_0_0_595 (.ZN (n_0_0_498), .A1 (n_0_0_497), .A2 (hfn_ipo_n63), .B1 (hfn_ipo_n81), .B2 (n_0_0_476));
OAI22_X1 i_0_0_594 (.ZN (n_0_0_497), .A1 (n_0_0_496), .A2 (hfn_ipo_n78), .B1 (n_0_0_450), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_593 (.ZN (n_0_0_496), .A1 (n_0_0_495), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_382));
AOI221_X1 i_0_0_592 (.ZN (n_0_0_495), .A (n_0_0_426), .B1 (\extended_M[20] ), .B2 (n_0_0_412)
    , .C1 (\extended_M[4] ), .C2 (n_0_0_442));
AOI22_X1 i_0_0_591 (.ZN (n_0_0_494), .A1 (hfn_ipo_n65), .A2 (n_0_0_493), .B1 (hfn_ipo_n69), .B2 (n_0_0_488));
OAI22_X1 i_0_0_590 (.ZN (n_0_0_493), .A1 (n_0_0_492), .A2 (hfn_ipo_n81), .B1 (n_0_0_470), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_589 (.ZN (n_0_0_492), .A1 (n_0_0_491), .A2 (hfn_ipo_n78), .B1 (n_0_0_445), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_588 (.ZN (n_0_0_491), .A1 (n_0_0_490), .A2 (hfn_ipo_n75), .B1 (n_0_0_8), .B2 (n_0_0_391));
AOI221_X1 i_0_0_587 (.ZN (n_0_0_490), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[4] )
    , .B2 (n_0_0_442), .C1 (\extended_M_mul_neg_one[20] ), .C2 (n_0_0_412));
NAND2_X1 i_0_0_586 (.ZN (\partialProd[35] ), .A1 (n_0_0_484), .A2 (n_0_0_489));
AOI22_X1 i_0_0_585 (.ZN (n_0_0_489), .A1 (hfn_ipo_n65), .A2 (n_0_0_488), .B1 (hfn_ipo_n69), .B2 (n_0_0_471));
AOI22_X1 i_0_0_584 (.ZN (n_0_0_488), .A1 (n_0_0_487), .A2 (hfn_ipo_n63), .B1 (n_0_0_457), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_583 (.ZN (n_0_0_487), .A1 (n_0_0_486), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_437));
OAI22_X1 i_0_0_582 (.ZN (n_0_0_486), .A1 (n_0_0_485), .A2 (hfn_ipo_n75), .B1 (n_0_0_8), .B2 (n_0_0_368));
AOI221_X1 i_0_0_581 (.ZN (n_0_0_485), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[3] )
    , .B2 (n_0_0_442), .C1 (\extended_M_mul_neg_one[19] ), .C2 (n_0_0_412));
AOI22_X1 i_0_0_580 (.ZN (n_0_0_484), .A1 (n_0_0_74), .A2 (n_0_0_483), .B1 (n_0_0_94), .B2 (n_0_0_477));
AOI22_X1 i_0_0_579 (.ZN (n_0_0_483), .A1 (n_0_0_482), .A2 (hfn_ipo_n63), .B1 (n_0_0_465), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_578 (.ZN (n_0_0_482), .A1 (n_0_0_481), .A2 (hfn_ipo_n78), .B1 (n_0_0_429), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_577 (.ZN (n_0_0_481), .A1 (n_0_0_480), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_376));
AOI22_X1 i_0_0_576 (.ZN (n_0_0_480), .A1 (n_0_0_461), .A2 (n_0_0_479), .B1 (\extended_M[19] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_575 (.ZN (n_0_0_479), .A1 (n_0_0_101), .A2 (drc_ipo_n84));
NAND2_X1 i_0_0_574 (.ZN (\partialProd[34] ), .A1 (n_0_0_472), .A2 (n_0_0_478));
AOI22_X1 i_0_0_573 (.ZN (n_0_0_478), .A1 (n_0_0_74), .A2 (n_0_0_477), .B1 (n_0_0_90), .B2 (n_0_0_458));
AOI22_X1 i_0_0_572 (.ZN (n_0_0_477), .A1 (n_0_0_451), .A2 (hfn_ipo_n81), .B1 (hfn_ipo_n63), .B2 (n_0_0_476));
OAI22_X1 i_0_0_571 (.ZN (n_0_0_476), .A1 (n_0_0_475), .A2 (hfn_ipo_n78), .B1 (n_0_0_421), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_570 (.ZN (n_0_0_475), .A1 (n_0_0_474), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_362));
AOI22_X1 i_0_0_569 (.ZN (n_0_0_474), .A1 (n_0_0_461), .A2 (n_0_0_473), .B1 (\extended_M[18] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_568 (.ZN (n_0_0_473), .A1 (n_0_0_107), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_567 (.ZN (n_0_0_472), .A1 (hfn_ipo_n65), .A2 (n_0_0_471), .B1 (n_0_0_94), .B2 (n_0_0_466));
AOI22_X1 i_0_0_566 (.ZN (n_0_0_471), .A1 (n_0_0_470), .A2 (hfn_ipo_n63), .B1 (n_0_0_446), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_565 (.ZN (n_0_0_470), .A1 (n_0_0_469), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_414));
OAI22_X1 i_0_0_564 (.ZN (n_0_0_469), .A1 (n_0_0_468), .A2 (hfn_ipo_n75), .B1 (n_0_0_8), .B2 (n_0_0_351));
AOI221_X1 i_0_0_563 (.ZN (n_0_0_468), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[2] )
    , .B2 (n_0_0_442), .C1 (\extended_M_mul_neg_one[18] ), .C2 (n_0_0_412));
NAND2_X1 i_0_0_562 (.ZN (\partialProd[33] ), .A1 (n_0_0_459), .A2 (n_0_0_467));
AOI22_X1 i_0_0_561 (.ZN (n_0_0_467), .A1 (n_0_0_74), .A2 (n_0_0_466), .B1 (n_0_0_90), .B2 (n_0_0_447));
AOI22_X1 i_0_0_560 (.ZN (n_0_0_466), .A1 (n_0_0_430), .A2 (hfn_ipo_n81), .B1 (n_0_0_465), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_559 (.ZN (n_0_0_465), .A1 (n_0_0_464), .A2 (hfn_ipo_n78), .B1 (n_0_0_407), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_558 (.ZN (n_0_0_464), .A1 (n_0_0_463), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_345));
AOI22_X1 i_0_0_557 (.ZN (n_0_0_463), .A1 (n_0_0_461), .A2 (n_0_0_462), .B1 (\extended_M[17] ), .B2 (n_0_0_412));
NAND2_X1 i_0_0_556 (.ZN (n_0_0_462), .A1 (n_0_0_147), .A2 (drc_ipo_n84));
NOR2_X1 i_0_0_555 (.ZN (n_0_0_461), .A1 (n_0_0_460), .A2 (drc_ipo_n83));
NOR2_X1 i_0_0_554 (.ZN (n_0_0_460), .A1 (\extended_M[63] ), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_553 (.ZN (n_0_0_459), .A1 (hfn_ipo_n65), .A2 (n_0_0_458), .B1 (n_0_0_94), .B2 (n_0_0_453));
AOI22_X1 i_0_0_552 (.ZN (n_0_0_458), .A1 (n_0_0_457), .A2 (hfn_ipo_n63), .B1 (hfn_ipo_n81), .B2 (n_0_0_438));
OAI22_X1 i_0_0_551 (.ZN (n_0_0_457), .A1 (n_0_0_456), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_401));
OAI22_X1 i_0_0_550 (.ZN (n_0_0_456), .A1 (n_0_0_455), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_336));
AOI221_X1 i_0_0_549 (.ZN (n_0_0_455), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[1] )
    , .B2 (n_0_0_442), .C1 (\extended_M_mul_neg_one[17] ), .C2 (n_0_0_412));
NAND2_X1 i_0_0_548 (.ZN (\partialProd[32] ), .A1 (n_0_0_448), .A2 (n_0_0_454));
AOI22_X1 i_0_0_547 (.ZN (n_0_0_454), .A1 (n_0_0_74), .A2 (n_0_0_453), .B1 (n_0_0_90), .B2 (n_0_0_439));
AOI22_X1 i_0_0_546 (.ZN (n_0_0_453), .A1 (n_0_0_451), .A2 (hfn_ipo_n63), .B1 (hfn_ipo_n81), .B2 (n_0_0_452));
INV_X1 i_0_0_545 (.ZN (n_0_0_452), .A (n_0_0_423));
OAI22_X1 i_0_0_544 (.ZN (n_0_0_451), .A1 (n_0_0_450), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_385));
OAI22_X1 i_0_0_543 (.ZN (n_0_0_450), .A1 (n_0_0_449), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_327));
AOI211_X1 i_0_0_542 (.ZN (n_0_0_449), .A (n_0_0_426), .B (n_0_0_443), .C1 (\extended_M[16] ), .C2 (n_0_0_412));
AOI22_X1 i_0_0_541 (.ZN (n_0_0_448), .A1 (hfn_ipo_n66), .A2 (n_0_0_447), .B1 (n_0_0_94), .B2 (n_0_0_432));
AOI22_X1 i_0_0_540 (.ZN (n_0_0_447), .A1 (n_0_0_446), .A2 (hfn_ipo_n63), .B1 (hfn_ipo_n81), .B2 (n_0_0_415));
OAI22_X1 i_0_0_539 (.ZN (n_0_0_446), .A1 (n_0_0_445), .A2 (hfn_ipo_n78), .B1 (hfn_ipo_n60), .B2 (n_0_0_394));
OAI22_X1 i_0_0_538 (.ZN (n_0_0_445), .A1 (n_0_0_444), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_322));
AOI211_X1 i_0_0_537 (.ZN (n_0_0_444), .A (n_0_0_435), .B (n_0_0_443), .C1 (\extended_M_mul_neg_one[16] ), .C2 (n_0_0_412));
AND2_X1 i_0_0_536 (.ZN (n_0_0_443), .A1 (n_0_0_442), .A2 (\extended_M[0] ));
NOR2_X2 i_0_0_535 (.ZN (n_0_0_442), .A1 (n_0_0_7), .A2 (drc_ipo_n83));
NAND2_X1 i_0_0_534 (.ZN (\partialProd[31] ), .A1 (n_0_0_433), .A2 (n_0_0_441));
AOI22_X1 i_0_0_533 (.ZN (n_0_0_441), .A1 (hfn_ipo_n66), .A2 (n_0_0_439), .B1 (n_0_0_94), .B2 (n_0_0_440));
INV_X1 i_0_0_532 (.ZN (n_0_0_440), .A (n_0_0_424));
AOI22_X1 i_0_0_531 (.ZN (n_0_0_439), .A1 (n_0_0_438), .A2 (hfn_ipo_n63), .B1 (n_0_0_402), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_0_530 (.ZN (n_0_0_438), .A1 (n_0_0_437), .A2 (hfn_ipo_n60), .B1 (n_0_0_371), .B2 (hfn_ipo_n78));
OAI22_X1 i_0_0_529 (.ZN (n_0_0_437), .A1 (n_0_0_436), .A2 (hfn_ipo_n76), .B1 (n_0_0_8), .B2 (n_0_0_311));
AOI21_X1 i_0_0_528 (.ZN (n_0_0_436), .A (n_0_0_435), .B1 (\extended_M_mul_neg_one[15] ), .B2 (n_0_0_412));
NOR2_X2 i_0_0_527 (.ZN (n_0_0_435), .A1 (n_0_0_434), .A2 (drc_ipo_n83));
NAND2_X1 i_0_0_526 (.ZN (n_0_0_434), .A1 (n_0_0_7), .A2 (\extended_M_mul_neg_one[63] ));
AOI22_X1 i_0_0_525 (.ZN (n_0_0_433), .A1 (n_0_0_74), .A2 (n_0_0_432), .B1 (n_0_0_90), .B2 (n_0_0_416));
AOI22_X1 i_0_0_524 (.ZN (n_0_0_432), .A1 (n_0_0_430), .A2 (hfn_ipo_n63), .B1 (n_0_0_431), .B2 (hfn_ipo_n81));
INV_X1 i_0_0_523 (.ZN (n_0_0_431), .A (n_0_0_409));
OAI22_X1 i_0_0_522 (.ZN (n_0_0_430), .A1 (n_0_0_429), .A2 (hfn_ipo_n78), .B1 (n_0_0_378), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_521 (.ZN (n_0_0_429), .A1 (n_0_0_427), .A2 (hfn_ipo_n76), .B1 (n_0_0_428), .B2 (n_0_0_318));
INV_X1 i_0_0_520 (.ZN (n_0_0_428), .A (n_0_0_317));
AOI21_X1 i_0_0_519 (.ZN (n_0_0_427), .A (n_0_0_426), .B1 (\extended_M[15] ), .B2 (n_0_0_412));
NOR2_X1 i_0_0_518 (.ZN (n_0_0_426), .A1 (n_0_0_425), .A2 (drc_ipo_n83));
NAND2_X1 i_0_0_517 (.ZN (n_0_0_425), .A1 (n_0_0_7), .A2 (\extended_M[63] ));
OAI221_X1 i_0_0_516 (.ZN (\partialProd[30] ), .A (n_0_0_417), .B1 (n_0_0_70), .B2 (n_0_0_410)
    , .C1 (n_0_0_73), .C2 (n_0_0_424));
OAI22_X1 i_0_0_515 (.ZN (n_0_0_424), .A1 (n_0_0_418), .A2 (hfn_ipo_n63), .B1 (n_0_0_423), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_0_514 (.ZN (n_0_0_423), .A1 (n_0_0_364), .A2 (hfn_ipo_n78), .B1 (n_0_0_422), .B2 (hfn_ipo_n60));
INV_X1 i_0_0_513 (.ZN (n_0_0_422), .A (n_0_0_421));
AND2_X1 i_0_0_512 (.ZN (n_0_0_421), .A1 (n_0_0_420), .A2 (n_0_0_7));
OAI22_X1 i_0_0_511 (.ZN (n_0_0_420), .A1 (n_0_0_305), .A2 (hfn_ipo_n73), .B1 (n_0_0_419), .B2 (hfn_ipo_n75));
AOI22_X1 i_0_0_510 (.ZN (n_0_0_419), .A1 (n_0_0_15), .A2 (\extended_M[30] ), .B1 (\extended_M[14] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_509 (.ZN (n_0_0_418), .A (n_0_0_386));
AOI22_X1 i_0_0_508 (.ZN (n_0_0_417), .A1 (hfn_ipo_n66), .A2 (n_0_0_416), .B1 (n_0_0_90), .B2 (n_0_0_403));
AOI22_X1 i_0_0_507 (.ZN (n_0_0_416), .A1 (n_0_0_415), .A2 (hfn_ipo_n63), .B1 (n_0_0_395), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_506 (.ZN (n_0_0_415), .A1 (n_0_0_414), .A2 (hfn_ipo_n78), .B1 (n_0_0_354), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_505 (.ZN (n_0_0_414), .A1 (n_0_0_300), .A2 (n_0_0_318), .B1 (n_0_0_413), .B2 (hfn_ipo_n76));
AOI22_X1 i_0_0_504 (.ZN (n_0_0_413), .A1 (n_0_0_411), .A2 (n_0_0_15), .B1 (n_0_0_412), .B2 (\extended_M_mul_neg_one[14] ));
NOR2_X4 i_0_0_503 (.ZN (n_0_0_412), .A1 (n_0_0_15), .A2 (drc_ipo_n84));
AND2_X1 i_0_0_502 (.ZN (n_0_0_411), .A1 (n_0_0_7), .A2 (\extended_M_mul_neg_one[30] ));
OAI221_X1 i_0_0_501 (.ZN (\partialProd[29] ), .A (n_0_0_404), .B1 (n_0_0_69), .B2 (n_0_0_397)
    , .C1 (n_0_0_73), .C2 (n_0_0_410));
AOI22_X1 i_0_0_500 (.ZN (n_0_0_410), .A1 (n_0_0_409), .A2 (hfn_ipo_n64), .B1 (n_0_0_380), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_0_499 (.ZN (n_0_0_409), .A1 (n_0_0_408), .A2 (hfn_ipo_n60), .B1 (n_0_0_347), .B2 (hfn_ipo_n79));
INV_X1 i_0_0_498 (.ZN (n_0_0_408), .A (n_0_0_407));
AND2_X1 i_0_0_497 (.ZN (n_0_0_407), .A1 (n_0_0_406), .A2 (n_0_0_7));
OAI22_X1 i_0_0_496 (.ZN (n_0_0_406), .A1 (n_0_0_318), .A2 (n_0_0_283), .B1 (n_0_0_405), .B2 (hfn_ipo_n76));
AOI22_X1 i_0_0_495 (.ZN (n_0_0_405), .A1 (n_0_0_15), .A2 (\extended_M[29] ), .B1 (\extended_M[13] ), .B2 (drc_ipo_n83));
AOI22_X1 i_0_0_494 (.ZN (n_0_0_404), .A1 (hfn_ipo_n66), .A2 (n_0_0_403), .B1 (n_0_0_94), .B2 (n_0_0_388));
AOI22_X1 i_0_0_493 (.ZN (n_0_0_403), .A1 (n_0_0_402), .A2 (hfn_ipo_n63), .B1 (n_0_0_372), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_492 (.ZN (n_0_0_402), .A1 (n_0_0_401), .A2 (hfn_ipo_n78), .B1 (n_0_0_339), .B2 (hfn_ipo_n60));
NOR2_X1 i_0_0_491 (.ZN (n_0_0_401), .A1 (n_0_0_400), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_490 (.ZN (n_0_0_400), .A1 (n_0_0_292), .A2 (hfn_ipo_n75), .B1 (n_0_0_399), .B2 (hfn_ipo_n73));
INV_X1 i_0_0_489 (.ZN (n_0_0_399), .A (n_0_0_398));
AOI22_X1 i_0_0_488 (.ZN (n_0_0_398), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[29] )
    , .B1 (\extended_M_mul_neg_one[13] ), .B2 (drc_ipo_n83));
OAI221_X1 i_0_0_487 (.ZN (\partialProd[28] ), .A (n_0_0_389), .B1 (n_0_0_70), .B2 (n_0_0_381)
    , .C1 (n_0_0_67), .C2 (n_0_0_397));
OAI22_X1 i_0_0_486 (.ZN (n_0_0_397), .A1 (n_0_0_396), .A2 (hfn_ipo_n81), .B1 (n_0_0_357), .B2 (hfn_ipo_n63));
INV_X1 i_0_0_485 (.ZN (n_0_0_396), .A (n_0_0_395));
OAI22_X1 i_0_0_484 (.ZN (n_0_0_395), .A1 (n_0_0_394), .A2 (hfn_ipo_n78), .B1 (n_0_0_323), .B2 (hfn_ipo_n60));
NOR2_X1 i_0_0_483 (.ZN (n_0_0_394), .A1 (n_0_0_393), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_482 (.ZN (n_0_0_393), .A1 (n_0_0_390), .A2 (hfn_ipo_n75), .B1 (n_0_0_392), .B2 (hfn_ipo_n73));
INV_X1 i_0_0_481 (.ZN (n_0_0_392), .A (n_0_0_391));
AOI22_X1 i_0_0_480 (.ZN (n_0_0_391), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[28] )
    , .B1 (\extended_M_mul_neg_one[12] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_479 (.ZN (n_0_0_390), .A (n_0_0_271));
AOI22_X1 i_0_0_478 (.ZN (n_0_0_389), .A1 (n_0_0_74), .A2 (n_0_0_388), .B1 (n_0_0_90), .B2 (n_0_0_373));
OAI22_X1 i_0_0_477 (.ZN (n_0_0_388), .A1 (n_0_0_386), .A2 (hfn_ipo_n81), .B1 (n_0_0_387), .B2 (hfn_ipo_n63));
INV_X1 i_0_0_476 (.ZN (n_0_0_387), .A (n_0_0_365));
OAI22_X1 i_0_0_475 (.ZN (n_0_0_386), .A1 (n_0_0_330), .A2 (hfn_ipo_n60), .B1 (n_0_0_385), .B2 (hfn_ipo_n78));
NOR2_X1 i_0_0_474 (.ZN (n_0_0_385), .A1 (n_0_0_384), .A2 (drc_ipo_n84));
OAI22_X1 i_0_0_473 (.ZN (n_0_0_384), .A1 (n_0_0_278), .A2 (n_0_0_318), .B1 (n_0_0_383), .B2 (hfn_ipo_n76));
INV_X1 i_0_0_472 (.ZN (n_0_0_383), .A (n_0_0_382));
AOI22_X1 i_0_0_471 (.ZN (n_0_0_382), .A1 (n_0_0_15), .A2 (\extended_M[28] ), .B1 (\extended_M[12] ), .B2 (drc_ipo_n83));
OAI21_X1 i_0_0_470 (.ZN (\partialProd[27] ), .A (n_0_0_375), .B1 (n_0_0_73), .B2 (n_0_0_381));
AOI22_X1 i_0_0_469 (.ZN (n_0_0_381), .A1 (n_0_0_380), .A2 (hfn_ipo_n64), .B1 (n_0_0_348), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_0_468 (.ZN (n_0_0_380), .A1 (n_0_0_379), .A2 (hfn_ipo_n61), .B1 (n_0_0_319), .B2 (hfn_ipo_n79));
INV_X1 i_0_0_467 (.ZN (n_0_0_379), .A (n_0_0_378));
AND2_X1 i_0_0_466 (.ZN (n_0_0_378), .A1 (n_0_0_377), .A2 (n_0_0_7));
AOI22_X1 i_0_0_465 (.ZN (n_0_0_377), .A1 (n_0_0_264), .A2 (hfn_ipo_n76), .B1 (n_0_0_376), .B2 (n_0_0_318));
AOI22_X1 i_0_0_464 (.ZN (n_0_0_376), .A1 (n_0_0_15), .A2 (\extended_M[27] ), .B1 (\extended_M[11] ), .B2 (drc_ipo_n83));
AOI222_X1 i_0_0_463 (.ZN (n_0_0_375), .A1 (hfn_ipo_n66), .A2 (n_0_0_373), .B1 (n_0_0_90)
    , .B2 (n_0_0_359), .C1 (n_0_0_94), .C2 (n_0_0_374));
INV_X1 i_0_0_462 (.ZN (n_0_0_374), .A (n_0_0_366));
OAI22_X1 i_0_0_461 (.ZN (n_0_0_373), .A1 (n_0_0_341), .A2 (hfn_ipo_n63), .B1 (n_0_0_372), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_0_460 (.ZN (n_0_0_372), .A1 (n_0_0_371), .A2 (hfn_ipo_n60), .B1 (n_0_0_312), .B2 (hfn_ipo_n78));
NOR2_X1 i_0_0_459 (.ZN (n_0_0_371), .A1 (n_0_0_370), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_458 (.ZN (n_0_0_370), .A1 (n_0_0_367), .A2 (hfn_ipo_n75), .B1 (n_0_0_369), .B2 (hfn_ipo_n73));
INV_X1 i_0_0_457 (.ZN (n_0_0_369), .A (n_0_0_368));
AOI22_X1 i_0_0_456 (.ZN (n_0_0_368), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[27] )
    , .B1 (\extended_M_mul_neg_one[11] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_455 (.ZN (n_0_0_367), .A (n_0_0_259));
OAI221_X1 i_0_0_454 (.ZN (\partialProd[26] ), .A (n_0_0_360), .B1 (n_0_0_70), .B2 (n_0_0_349)
    , .C1 (n_0_0_73), .C2 (n_0_0_366));
OAI22_X1 i_0_0_453 (.ZN (n_0_0_366), .A1 (n_0_0_361), .A2 (hfn_ipo_n64), .B1 (n_0_0_365), .B2 (hfn_ipo_n81));
AOI22_X1 i_0_0_452 (.ZN (n_0_0_365), .A1 (n_0_0_364), .A2 (hfn_ipo_n61), .B1 (n_0_0_307), .B2 (hfn_ipo_n79));
NAND2_X1 i_0_0_451 (.ZN (n_0_0_364), .A1 (n_0_0_363), .A2 (n_0_0_7));
OAI22_X1 i_0_0_450 (.ZN (n_0_0_363), .A1 (n_0_0_247), .A2 (n_0_0_318), .B1 (n_0_0_362), .B2 (hfn_ipo_n76));
AOI22_X1 i_0_0_449 (.ZN (n_0_0_362), .A1 (n_0_0_15), .A2 (\extended_M[26] ), .B1 (\extended_M[10] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_448 (.ZN (n_0_0_361), .A (n_0_0_332));
AOI22_X1 i_0_0_447 (.ZN (n_0_0_360), .A1 (hfn_ipo_n66), .A2 (n_0_0_359), .B1 (n_0_0_90), .B2 (n_0_0_342));
OAI22_X1 i_0_0_446 (.ZN (n_0_0_359), .A1 (n_0_0_358), .A2 (hfn_ipo_n82), .B1 (n_0_0_324), .B2 (hfn_ipo_n64));
INV_X1 i_0_0_445 (.ZN (n_0_0_358), .A (n_0_0_357));
OAI22_X1 i_0_0_444 (.ZN (n_0_0_357), .A1 (n_0_0_355), .A2 (hfn_ipo_n79), .B1 (n_0_0_356), .B2 (hfn_ipo_n60));
INV_X1 i_0_0_443 (.ZN (n_0_0_356), .A (n_0_0_301));
INV_X1 i_0_0_442 (.ZN (n_0_0_355), .A (n_0_0_354));
NOR2_X1 i_0_0_441 (.ZN (n_0_0_354), .A1 (n_0_0_353), .A2 (drc_ipo_n84));
AOI22_X1 i_0_0_440 (.ZN (n_0_0_353), .A1 (n_0_0_350), .A2 (hfn_ipo_n75), .B1 (n_0_0_352), .B2 (hfn_ipo_n73));
INV_X1 i_0_0_439 (.ZN (n_0_0_352), .A (n_0_0_351));
AOI22_X1 i_0_0_438 (.ZN (n_0_0_351), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[26] )
    , .B1 (\extended_M_mul_neg_one[10] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_437 (.ZN (n_0_0_350), .A (n_0_0_254));
OAI221_X1 i_0_0_436 (.ZN (\partialProd[25] ), .A (n_0_0_343), .B1 (n_0_0_69), .B2 (n_0_0_344)
    , .C1 (n_0_0_73), .C2 (n_0_0_349));
AOI22_X1 i_0_0_435 (.ZN (n_0_0_349), .A1 (n_0_0_320), .A2 (hfn_ipo_n82), .B1 (n_0_0_348), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_434 (.ZN (n_0_0_348), .A1 (n_0_0_347), .A2 (hfn_ipo_n79), .B1 (n_0_0_285), .B2 (hfn_ipo_n60));
AOI22_X1 i_0_0_433 (.ZN (n_0_0_347), .A1 (n_0_0_241), .A2 (hfn_ipo_n76), .B1 (n_0_0_346), .B2 (n_0_0_10));
INV_X1 i_0_0_432 (.ZN (n_0_0_346), .A (n_0_0_345));
OAI22_X1 i_0_0_431 (.ZN (n_0_0_345), .A1 (n_0_0_15), .A2 (\extended_M[9] ), .B1 (\extended_M[25] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_430 (.ZN (n_0_0_344), .A (n_0_0_325));
AOI22_X1 i_0_0_429 (.ZN (n_0_0_343), .A1 (hfn_ipo_n66), .A2 (n_0_0_342), .B1 (n_0_0_94), .B2 (n_0_0_334));
AOI22_X1 i_0_0_428 (.ZN (n_0_0_342), .A1 (n_0_0_341), .A2 (hfn_ipo_n63), .B1 (n_0_0_313), .B2 (hfn_ipo_n81));
OAI22_X1 i_0_0_427 (.ZN (n_0_0_341), .A1 (n_0_0_339), .A2 (hfn_ipo_n78), .B1 (n_0_0_340), .B2 (hfn_ipo_n60));
INV_X1 i_0_0_426 (.ZN (n_0_0_340), .A (n_0_0_293));
NOR2_X1 i_0_0_425 (.ZN (n_0_0_339), .A1 (n_0_0_338), .A2 (drc_ipo_n84));
OAI22_X1 i_0_0_424 (.ZN (n_0_0_338), .A1 (n_0_0_234), .A2 (n_0_0_318), .B1 (n_0_0_337), .B2 (hfn_ipo_n76));
INV_X1 i_0_0_423 (.ZN (n_0_0_337), .A (n_0_0_336));
AOI22_X1 i_0_0_422 (.ZN (n_0_0_336), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[25] )
    , .B1 (\extended_M_mul_neg_one[9] ), .B2 (drc_ipo_n83));
OAI221_X1 i_0_0_421 (.ZN (\partialProd[24] ), .A (n_0_0_326), .B1 (n_0_0_70), .B2 (n_0_0_321)
    , .C1 (n_0_0_73), .C2 (n_0_0_335));
INV_X1 i_0_0_420 (.ZN (n_0_0_335), .A (n_0_0_334));
OAI22_X1 i_0_0_419 (.ZN (n_0_0_334), .A1 (n_0_0_332), .A2 (hfn_ipo_n81), .B1 (n_0_0_333), .B2 (hfn_ipo_n63));
INV_X1 i_0_0_418 (.ZN (n_0_0_333), .A (n_0_0_308));
AOI22_X1 i_0_0_417 (.ZN (n_0_0_332), .A1 (n_0_0_330), .A2 (hfn_ipo_n60), .B1 (n_0_0_331), .B2 (hfn_ipo_n79));
INV_X1 i_0_0_416 (.ZN (n_0_0_331), .A (n_0_0_279));
NOR2_X1 i_0_0_415 (.ZN (n_0_0_330), .A1 (n_0_0_329), .A2 (drc_ipo_n84));
OAI22_X1 i_0_0_414 (.ZN (n_0_0_329), .A1 (n_0_0_220), .A2 (n_0_0_318), .B1 (n_0_0_328), .B2 (hfn_ipo_n76));
INV_X1 i_0_0_413 (.ZN (n_0_0_328), .A (n_0_0_327));
AOI22_X1 i_0_0_412 (.ZN (n_0_0_327), .A1 (n_0_0_15), .A2 (\extended_M[24] ), .B1 (\extended_M[8] ), .B2 (drc_ipo_n83));
AOI22_X1 i_0_0_411 (.ZN (n_0_0_326), .A1 (hfn_ipo_n66), .A2 (n_0_0_325), .B1 (n_0_0_90), .B2 (n_0_0_314));
AOI22_X1 i_0_0_410 (.ZN (n_0_0_325), .A1 (n_0_0_302), .A2 (hfn_ipo_n82), .B1 (n_0_0_324), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_409 (.ZN (n_0_0_324), .A1 (n_0_0_323), .A2 (hfn_ipo_n78), .B1 (n_0_0_272), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_408 (.ZN (n_0_0_323), .A1 (n_0_0_228), .A2 (n_0_0_318), .B1 (n_0_0_322), .B2 (n_0_0_14));
AOI22_X1 i_0_0_407 (.ZN (n_0_0_322), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[24] )
    , .B1 (\extended_M_mul_neg_one[8] ), .B2 (drc_ipo_n83));
OAI221_X1 i_0_0_406 (.ZN (\partialProd[23] ), .A (n_0_0_315), .B1 (n_0_0_70), .B2 (n_0_0_309)
    , .C1 (n_0_0_73), .C2 (n_0_0_321));
AOI22_X1 i_0_0_405 (.ZN (n_0_0_321), .A1 (n_0_0_320), .A2 (hfn_ipo_n64), .B1 (n_0_0_286), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_0_404 (.ZN (n_0_0_320), .A1 (n_0_0_319), .A2 (hfn_ipo_n61), .B1 (n_0_0_266), .B2 (hfn_ipo_n79));
AOI22_X1 i_0_0_403 (.ZN (n_0_0_319), .A1 (n_0_0_317), .A2 (n_0_0_318), .B1 (n_0_0_128), .B2 (\extended_M[15] ));
INV_X1 i_0_0_402 (.ZN (n_0_0_318), .A (hfn_ipo_n75));
NOR2_X1 i_0_0_401 (.ZN (n_0_0_317), .A1 (n_0_0_316), .A2 (drc_ipo_n84));
OAI22_X1 i_0_0_400 (.ZN (n_0_0_316), .A1 (n_0_0_15), .A2 (\extended_M[7] ), .B1 (\extended_M[23] ), .B2 (drc_ipo_n83));
AOI22_X1 i_0_0_399 (.ZN (n_0_0_315), .A1 (hfn_ipo_n66), .A2 (n_0_0_314), .B1 (n_0_0_90), .B2 (n_0_0_303));
AOI22_X1 i_0_0_398 (.ZN (n_0_0_314), .A1 (hfn_ipo_n81), .A2 (n_0_0_310), .B1 (n_0_0_313), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_397 (.ZN (n_0_0_313), .A1 (n_0_0_312), .A2 (hfn_ipo_n79), .B1 (n_0_0_260), .B2 (hfn_ipo_n60));
OAI22_X1 i_0_0_396 (.ZN (n_0_0_312), .A1 (n_0_0_140), .A2 (n_0_0_208), .B1 (n_0_0_311), .B2 (n_0_0_14));
AOI22_X1 i_0_0_395 (.ZN (n_0_0_311), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[23] )
    , .B1 (\extended_M_mul_neg_one[7] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_394 (.ZN (n_0_0_310), .A (n_0_0_294));
OAI221_X1 i_0_0_393 (.ZN (\partialProd[22] ), .A (n_0_0_297), .B1 (n_0_0_67), .B2 (n_0_0_304)
    , .C1 (n_0_0_73), .C2 (n_0_0_309));
AOI22_X1 i_0_0_392 (.ZN (n_0_0_309), .A1 (n_0_0_280), .A2 (hfn_ipo_n81), .B1 (n_0_0_308), .B2 (hfn_ipo_n63));
OAI22_X1 i_0_0_391 (.ZN (n_0_0_308), .A1 (n_0_0_249), .A2 (hfn_ipo_n61), .B1 (n_0_0_307), .B2 (hfn_ipo_n79));
AOI22_X1 i_0_0_390 (.ZN (n_0_0_307), .A1 (n_0_0_306), .A2 (n_0_0_10), .B1 (n_0_0_128), .B2 (\extended_M[14] ));
INV_X1 i_0_0_389 (.ZN (n_0_0_306), .A (n_0_0_305));
OAI22_X1 i_0_0_388 (.ZN (n_0_0_305), .A1 (n_0_0_15), .A2 (\extended_M[6] ), .B1 (\extended_M[22] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_387 (.ZN (n_0_0_304), .A (n_0_0_303));
AOI22_X1 i_0_0_386 (.ZN (n_0_0_303), .A1 (n_0_0_302), .A2 (hfn_ipo_n64), .B1 (n_0_0_273), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_0_385 (.ZN (n_0_0_302), .A1 (n_0_0_301), .A2 (hfn_ipo_n61), .B1 (n_0_0_255), .B2 (hfn_ipo_n79));
OAI22_X1 i_0_0_384 (.ZN (n_0_0_301), .A1 (n_0_0_300), .A2 (hfn_ipo_n76), .B1 (n_0_0_140), .B2 (n_0_0_197));
NAND2_X1 i_0_0_383 (.ZN (n_0_0_300), .A1 (n_0_0_299), .A2 (n_0_0_7));
OAI22_X1 i_0_0_382 (.ZN (n_0_0_299), .A1 (n_0_0_115), .A2 (n_0_0_15), .B1 (n_0_0_298), .B2 (drc_ipo_n83));
INV_X1 i_0_0_381 (.ZN (n_0_0_298), .A (\extended_M_mul_neg_one[22] ));
AOI22_X1 i_0_0_380 (.ZN (n_0_0_297), .A1 (n_0_0_94), .A2 (n_0_0_288), .B1 (n_0_0_90), .B2 (n_0_0_296));
INV_X1 i_0_0_379 (.ZN (n_0_0_296), .A (n_0_0_295));
OAI221_X1 i_0_0_378 (.ZN (\partialProd[21] ), .A (n_0_0_289), .B1 (n_0_0_70), .B2 (n_0_0_281)
    , .C1 (n_0_0_67), .C2 (n_0_0_295));
OAI22_X1 i_0_0_377 (.ZN (n_0_0_295), .A1 (n_0_0_290), .A2 (hfn_ipo_n64), .B1 (n_0_0_294), .B2 (hfn_ipo_n82));
OAI22_X1 i_0_0_376 (.ZN (n_0_0_294), .A1 (n_0_0_293), .A2 (hfn_ipo_n79), .B1 (n_0_0_235), .B2 (hfn_ipo_n60));
AOI22_X1 i_0_0_375 (.ZN (n_0_0_293), .A1 (n_0_0_292), .A2 (n_0_0_10), .B1 (n_0_0_128), .B2 (\extended_M_mul_neg_one[13] ));
AOI22_X1 i_0_0_374 (.ZN (n_0_0_292), .A1 (n_0_0_291), .A2 (n_0_0_15), .B1 (n_0_0_191), .B2 (drc_ipo_n83));
INV_X1 i_0_0_373 (.ZN (n_0_0_291), .A (\extended_M_mul_neg_one[21] ));
INV_X1 i_0_0_372 (.ZN (n_0_0_290), .A (n_0_0_261));
AOI22_X1 i_0_0_371 (.ZN (n_0_0_289), .A1 (n_0_0_74), .A2 (n_0_0_288), .B1 (n_0_0_90), .B2 (n_0_0_274));
OAI22_X1 i_0_0_370 (.ZN (n_0_0_288), .A1 (n_0_0_287), .A2 (hfn_ipo_n82), .B1 (n_0_0_268), .B2 (hfn_ipo_n64));
INV_X1 i_0_0_369 (.ZN (n_0_0_287), .A (n_0_0_286));
OAI22_X1 i_0_0_368 (.ZN (n_0_0_286), .A1 (n_0_0_282), .A2 (hfn_ipo_n61), .B1 (n_0_0_285), .B2 (hfn_ipo_n79));
AOI22_X1 i_0_0_367 (.ZN (n_0_0_285), .A1 (n_0_0_10), .A2 (n_0_0_284), .B1 (n_0_0_128), .B2 (\extended_M[13] ));
INV_X1 i_0_0_366 (.ZN (n_0_0_284), .A (n_0_0_283));
OAI22_X1 i_0_0_365 (.ZN (n_0_0_283), .A1 (n_0_0_15), .A2 (\extended_M[5] ), .B1 (\extended_M[21] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_364 (.ZN (n_0_0_282), .A (n_0_0_243));
OAI221_X1 i_0_0_363 (.ZN (\partialProd[20] ), .A (n_0_0_275), .B1 (n_0_0_69), .B2 (n_0_0_276)
    , .C1 (n_0_0_73), .C2 (n_0_0_281));
AOI22_X1 i_0_0_362 (.ZN (n_0_0_281), .A1 (n_0_0_280), .A2 (hfn_ipo_n64), .B1 (n_0_0_250), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_0_361 (.ZN (n_0_0_280), .A1 (n_0_0_221), .A2 (hfn_ipo_n79), .B1 (n_0_0_279), .B2 (hfn_ipo_n60));
AOI22_X1 i_0_0_360 (.ZN (n_0_0_279), .A1 (n_0_0_278), .A2 (n_0_0_10), .B1 (n_0_0_128), .B2 (\extended_M[12] ));
INV_X1 i_0_0_359 (.ZN (n_0_0_278), .A (n_0_0_277));
AOI22_X1 i_0_0_358 (.ZN (n_0_0_277), .A1 (n_0_0_15), .A2 (\extended_M[20] ), .B1 (\extended_M[4] ), .B2 (drc_ipo_n83));
INV_X1 i_0_0_357 (.ZN (n_0_0_276), .A (n_0_0_262));
AOI22_X1 i_0_0_356 (.ZN (n_0_0_275), .A1 (hfn_ipo_n66), .A2 (n_0_0_274), .B1 (n_0_0_94), .B2 (n_0_0_269));
AOI22_X1 i_0_0_355 (.ZN (n_0_0_274), .A1 (n_0_0_273), .A2 (hfn_ipo_n64), .B1 (n_0_0_256), .B2 (hfn_ipo_n82));
OAI22_X1 i_0_0_354 (.ZN (n_0_0_273), .A1 (n_0_0_229), .A2 (hfn_ipo_n61), .B1 (n_0_0_272), .B2 (hfn_ipo_n79));
OAI22_X1 i_0_0_353 (.ZN (n_0_0_272), .A1 (n_0_0_140), .A2 (n_0_0_174), .B1 (n_0_0_271), .B2 (n_0_0_14));
OAI22_X1 i_0_0_352 (.ZN (n_0_0_271), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[4] )
    , .B1 (\extended_M_mul_neg_one[20] ), .B2 (drc_ipo_n83));
NAND2_X1 i_0_0_351 (.ZN (\partialProd[19] ), .A1 (n_0_0_263), .A2 (n_0_0_270));
AOI22_X1 i_0_0_350 (.ZN (n_0_0_270), .A1 (n_0_0_74), .A2 (n_0_0_269), .B1 (n_0_0_90), .B2 (n_0_0_257));
AOI22_X1 i_0_0_349 (.ZN (n_0_0_269), .A1 (n_0_0_244), .A2 (hfn_ipo_n82), .B1 (n_0_0_268), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_348 (.ZN (n_0_0_268), .A1 (n_0_0_267), .A2 (hfn_ipo_n79), .B1 (n_0_0_214), .B2 (hfn_ipo_n61));
INV_X1 i_0_0_347 (.ZN (n_0_0_267), .A (n_0_0_266));
AOI22_X1 i_0_0_346 (.ZN (n_0_0_266), .A1 (n_0_0_265), .A2 (n_0_0_10), .B1 (n_0_0_128), .B2 (\extended_M[11] ));
INV_X1 i_0_0_345 (.ZN (n_0_0_265), .A (n_0_0_264));
OAI22_X1 i_0_0_344 (.ZN (n_0_0_264), .A1 (n_0_0_15), .A2 (\extended_M[3] ), .B1 (\extended_M[19] ), .B2 (drc_ipo_n83));
AOI22_X1 i_0_0_343 (.ZN (n_0_0_263), .A1 (hfn_ipo_n66), .A2 (n_0_0_262), .B1 (n_0_0_94), .B2 (n_0_0_252));
AOI22_X1 i_0_0_342 (.ZN (n_0_0_262), .A1 (n_0_0_261), .A2 (hfn_ipo_n64), .B1 (n_0_0_237), .B2 (hfn_ipo_n82));
OAI22_X1 i_0_0_341 (.ZN (n_0_0_261), .A1 (n_0_0_260), .A2 (hfn_ipo_n79), .B1 (n_0_0_209), .B2 (hfn_ipo_n61));
OAI22_X1 i_0_0_340 (.ZN (n_0_0_260), .A1 (n_0_0_140), .A2 (n_0_0_168), .B1 (n_0_0_259), .B2 (n_0_0_14));
OAI22_X1 i_0_0_339 (.ZN (n_0_0_259), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[3] )
    , .B1 (\extended_M_mul_neg_one[19] ), .B2 (drc_ipo_n83));
NAND2_X1 i_0_0_338 (.ZN (\partialProd[18] ), .A1 (n_0_0_253), .A2 (n_0_0_258));
AOI22_X1 i_0_0_337 (.ZN (n_0_0_258), .A1 (hfn_ipo_n66), .A2 (n_0_0_257), .B1 (n_0_0_94), .B2 (n_0_0_245));
AOI22_X1 i_0_0_336 (.ZN (n_0_0_257), .A1 (n_0_0_230), .A2 (hfn_ipo_n82), .B1 (n_0_0_256), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_335 (.ZN (n_0_0_256), .A1 (n_0_0_255), .A2 (hfn_ipo_n79), .B1 (n_0_0_198), .B2 (hfn_ipo_n61));
OAI22_X1 i_0_0_334 (.ZN (n_0_0_255), .A1 (n_0_0_140), .A2 (n_0_0_158), .B1 (n_0_0_254), .B2 (n_0_0_14));
OAI22_X1 i_0_0_333 (.ZN (n_0_0_254), .A1 (n_0_0_15), .A2 (\extended_M_mul_neg_one[2] )
    , .B1 (\extended_M_mul_neg_one[18] ), .B2 (drc_ipo_n83));
AOI22_X1 i_0_0_332 (.ZN (n_0_0_253), .A1 (n_0_0_74), .A2 (n_0_0_252), .B1 (n_0_0_90), .B2 (n_0_0_238));
OAI22_X1 i_0_0_331 (.ZN (n_0_0_252), .A1 (n_0_0_223), .A2 (hfn_ipo_n64), .B1 (n_0_0_251), .B2 (hfn_ipo_n82));
INV_X1 i_0_0_330 (.ZN (n_0_0_251), .A (n_0_0_250));
OAI22_X1 i_0_0_329 (.ZN (n_0_0_250), .A1 (n_0_0_249), .A2 (hfn_ipo_n79), .B1 (n_0_0_202), .B2 (hfn_ipo_n61));
AOI22_X1 i_0_0_328 (.ZN (n_0_0_249), .A1 (n_0_0_10), .A2 (n_0_0_248), .B1 (n_0_0_128), .B2 (\extended_M[10] ));
INV_X1 i_0_0_327 (.ZN (n_0_0_248), .A (n_0_0_247));
OAI22_X1 i_0_0_326 (.ZN (n_0_0_247), .A1 (n_0_0_15), .A2 (\extended_M[2] ), .B1 (\extended_M[18] ), .B2 (drc_ipo_n83));
NAND2_X1 i_0_0_325 (.ZN (\partialProd[17] ), .A1 (n_0_0_239), .A2 (n_0_0_246));
AOI22_X1 i_0_0_324 (.ZN (n_0_0_246), .A1 (n_0_0_74), .A2 (n_0_0_245), .B1 (n_0_0_94), .B2 (n_0_0_224));
AOI22_X1 i_0_0_323 (.ZN (n_0_0_245), .A1 (n_0_0_244), .A2 (hfn_ipo_n64), .B1 (n_0_0_215), .B2 (hfn_ipo_n82));
OAI22_X1 i_0_0_322 (.ZN (n_0_0_244), .A1 (n_0_0_243), .A2 (hfn_ipo_n79), .B1 (n_0_0_187), .B2 (hfn_ipo_n61));
OAI22_X1 i_0_0_321 (.ZN (n_0_0_243), .A1 (n_0_0_242), .A2 (hfn_ipo_n76), .B1 (n_0_0_140), .B2 (n_0_0_148));
INV_X1 i_0_0_320 (.ZN (n_0_0_242), .A (n_0_0_241));
NOR2_X1 i_0_0_319 (.ZN (n_0_0_241), .A1 (n_0_0_240), .A2 (drc_ipo_n84));
OAI22_X1 i_0_0_318 (.ZN (n_0_0_240), .A1 (n_0_0_15), .A2 (\extended_M[1] ), .B1 (\extended_M[17] ), .B2 (drc_ipo_n83));
AOI22_X1 i_0_0_317 (.ZN (n_0_0_239), .A1 (hfn_ipo_n66), .A2 (n_0_0_238), .B1 (n_0_0_90), .B2 (n_0_0_231));
OAI22_X1 i_0_0_316 (.ZN (n_0_0_238), .A1 (n_0_0_237), .A2 (hfn_ipo_n82), .B1 (n_0_0_210), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_315 (.ZN (n_0_0_237), .A1 (n_0_0_236), .A2 (hfn_ipo_n79), .B1 (n_0_0_193), .B2 (hfn_ipo_n61));
INV_X1 i_0_0_314 (.ZN (n_0_0_236), .A (n_0_0_235));
AOI22_X1 i_0_0_313 (.ZN (n_0_0_235), .A1 (n_0_0_10), .A2 (n_0_0_234), .B1 (n_0_0_128), .B2 (\extended_M_mul_neg_one[9] ));
AOI22_X1 i_0_0_312 (.ZN (n_0_0_234), .A1 (n_0_0_233), .A2 (n_0_0_15), .B1 (n_0_0_141), .B2 (drc_ipo_n83));
INV_X1 i_0_0_311 (.ZN (n_0_0_233), .A (\extended_M_mul_neg_one[17] ));
NAND2_X1 i_0_0_310 (.ZN (\partialProd[16] ), .A1 (n_0_0_225), .A2 (n_0_0_232));
AOI22_X1 i_0_0_309 (.ZN (n_0_0_232), .A1 (hfn_ipo_n66), .A2 (n_0_0_231), .B1 (n_0_0_90), .B2 (n_0_0_211));
AOI22_X1 i_0_0_308 (.ZN (n_0_0_231), .A1 (n_0_0_230), .A2 (hfn_ipo_n64), .B1 (n_0_0_199), .B2 (hfn_ipo_n82));
OAI22_X1 i_0_0_307 (.ZN (n_0_0_230), .A1 (n_0_0_229), .A2 (hfn_ipo_n79), .B1 (n_0_0_175), .B2 (hfn_ipo_n61));
OAI22_X1 i_0_0_306 (.ZN (n_0_0_229), .A1 (n_0_0_228), .A2 (hfn_ipo_n76), .B1 (n_0_0_140), .B2 (n_0_0_130));
NAND2_X1 i_0_0_305 (.ZN (n_0_0_228), .A1 (n_0_0_227), .A2 (n_0_0_7));
OAI21_X1 i_0_0_304 (.ZN (n_0_0_227), .A (n_0_0_218), .B1 (n_0_0_226), .B2 (drc_ipo_n83));
INV_X1 i_0_0_303 (.ZN (n_0_0_226), .A (\extended_M_mul_neg_one[16] ));
AOI22_X1 i_0_0_302 (.ZN (n_0_0_225), .A1 (n_0_0_74), .A2 (n_0_0_224), .B1 (n_0_0_94), .B2 (n_0_0_216));
AOI22_X1 i_0_0_301 (.ZN (n_0_0_224), .A1 (n_0_0_223), .A2 (hfn_ipo_n64), .B1 (n_0_0_204), .B2 (hfn_ipo_n82));
OAI22_X1 i_0_0_300 (.ZN (n_0_0_223), .A1 (n_0_0_222), .A2 (hfn_ipo_n79), .B1 (n_0_0_181), .B2 (hfn_ipo_n61));
INV_X1 i_0_0_299 (.ZN (n_0_0_222), .A (n_0_0_221));
AOI22_X1 i_0_0_298 (.ZN (n_0_0_221), .A1 (n_0_0_220), .A2 (n_0_0_10), .B1 (n_0_0_128), .B2 (\extended_M[8] ));
OAI21_X1 i_0_0_297 (.ZN (n_0_0_220), .A (n_0_0_218), .B1 (n_0_0_219), .B2 (drc_ipo_n83));
INV_X1 i_0_0_296 (.ZN (n_0_0_219), .A (\extended_M[16] ));
NAND2_X1 i_0_0_295 (.ZN (n_0_0_218), .A1 (\extended_M[0] ), .A2 (drc_ipo_n83));
NAND2_X1 i_0_0_294 (.ZN (\partialProd[15] ), .A1 (n_0_0_212), .A2 (n_0_0_217));
AOI22_X1 i_0_0_293 (.ZN (n_0_0_217), .A1 (n_0_0_74), .A2 (n_0_0_216), .B1 (n_0_0_90), .B2 (n_0_0_200));
AOI22_X1 i_0_0_292 (.ZN (n_0_0_216), .A1 (n_0_0_188), .A2 (hfn_ipo_n82), .B1 (n_0_0_215), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_291 (.ZN (n_0_0_215), .A1 (n_0_0_214), .A2 (hfn_ipo_n79), .B1 (n_0_0_164), .B2 (hfn_ipo_n61));
OAI22_X1 i_0_0_290 (.ZN (n_0_0_214), .A1 (n_0_0_140), .A2 (n_0_0_120), .B1 (n_0_0_86), .B2 (n_0_0_213));
INV_X1 i_0_0_289 (.ZN (n_0_0_213), .A (\extended_M[15] ));
AOI22_X1 i_0_0_288 (.ZN (n_0_0_212), .A1 (hfn_ipo_n66), .A2 (n_0_0_211), .B1 (n_0_0_94), .B2 (n_0_0_205));
AOI22_X1 i_0_0_287 (.ZN (n_0_0_211), .A1 (hfn_ipo_n64), .A2 (n_0_0_210), .B1 (n_0_0_194), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_0_286 (.ZN (n_0_0_210), .A1 (n_0_0_209), .A2 (hfn_ipo_n61), .B1 (n_0_0_169), .B2 (hfn_ipo_n79));
OAI22_X1 i_0_0_285 (.ZN (n_0_0_209), .A1 (n_0_0_140), .A2 (n_0_0_207), .B1 (n_0_0_86), .B2 (n_0_0_208));
INV_X1 i_0_0_284 (.ZN (n_0_0_208), .A (\extended_M_mul_neg_one[15] ));
INV_X1 i_0_0_283 (.ZN (n_0_0_207), .A (\extended_M_mul_neg_one[7] ));
NAND2_X1 i_0_0_282 (.ZN (\partialProd[14] ), .A1 (n_0_0_201), .A2 (n_0_0_206));
AOI22_X1 i_0_0_281 (.ZN (n_0_0_206), .A1 (n_0_0_74), .A2 (n_0_0_205), .B1 (n_0_0_94), .B2 (n_0_0_189));
AOI22_X1 i_0_0_280 (.ZN (n_0_0_205), .A1 (n_0_0_182), .A2 (hfn_ipo_n82), .B1 (n_0_0_204), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_279 (.ZN (n_0_0_204), .A1 (n_0_0_203), .A2 (hfn_ipo_n79), .B1 (n_0_0_154), .B2 (hfn_ipo_n61));
INV_X1 i_0_0_278 (.ZN (n_0_0_203), .A (n_0_0_202));
AOI22_X1 i_0_0_277 (.ZN (n_0_0_202), .A1 (n_0_0_85), .A2 (\extended_M[14] ), .B1 (n_0_0_128), .B2 (\extended_M[6] ));
AOI22_X1 i_0_0_276 (.ZN (n_0_0_201), .A1 (hfn_ipo_n66), .A2 (n_0_0_200), .B1 (n_0_0_90), .B2 (n_0_0_195));
AOI22_X1 i_0_0_275 (.ZN (n_0_0_200), .A1 (n_0_0_176), .A2 (hfn_ipo_n82), .B1 (n_0_0_199), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_274 (.ZN (n_0_0_199), .A1 (n_0_0_198), .A2 (hfn_ipo_n79), .B1 (n_0_0_159), .B2 (hfn_ipo_n61));
OAI22_X1 i_0_0_273 (.ZN (n_0_0_198), .A1 (n_0_0_140), .A2 (n_0_0_115), .B1 (n_0_0_86), .B2 (n_0_0_197));
INV_X1 i_0_0_272 (.ZN (n_0_0_197), .A (\extended_M_mul_neg_one[14] ));
NAND2_X1 i_0_0_271 (.ZN (\partialProd[13] ), .A1 (n_0_0_190), .A2 (n_0_0_196));
AOI22_X1 i_0_0_270 (.ZN (n_0_0_196), .A1 (hfn_ipo_n66), .A2 (n_0_0_195), .B1 (n_0_0_90), .B2 (n_0_0_177));
OAI22_X1 i_0_0_269 (.ZN (n_0_0_195), .A1 (n_0_0_194), .A2 (hfn_ipo_n82), .B1 (n_0_0_170), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_268 (.ZN (n_0_0_194), .A1 (n_0_0_143), .A2 (hfn_ipo_n61), .B1 (n_0_0_193), .B2 (hfn_ipo_n79));
OAI22_X1 i_0_0_267 (.ZN (n_0_0_193), .A1 (n_0_0_140), .A2 (n_0_0_191), .B1 (n_0_0_86), .B2 (n_0_0_192));
INV_X1 i_0_0_266 (.ZN (n_0_0_192), .A (\extended_M_mul_neg_one[13] ));
INV_X1 i_0_0_265 (.ZN (n_0_0_191), .A (\extended_M_mul_neg_one[5] ));
AOI22_X1 i_0_0_264 (.ZN (n_0_0_190), .A1 (n_0_0_74), .A2 (n_0_0_189), .B1 (n_0_0_94), .B2 (n_0_0_183));
OAI22_X1 i_0_0_263 (.ZN (n_0_0_189), .A1 (n_0_0_188), .A2 (hfn_ipo_n82), .B1 (n_0_0_165), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_262 (.ZN (n_0_0_188), .A1 (n_0_0_149), .A2 (hfn_ipo_n61), .B1 (n_0_0_187), .B2 (hfn_ipo_n79));
OAI22_X1 i_0_0_261 (.ZN (n_0_0_187), .A1 (n_0_0_140), .A2 (n_0_0_185), .B1 (n_0_0_86), .B2 (n_0_0_186));
INV_X1 i_0_0_260 (.ZN (n_0_0_186), .A (\extended_M[13] ));
INV_X1 i_0_0_259 (.ZN (n_0_0_185), .A (\extended_M[5] ));
NAND2_X1 i_0_0_258 (.ZN (\partialProd[12] ), .A1 (n_0_0_178), .A2 (n_0_0_184));
AOI22_X1 i_0_0_257 (.ZN (n_0_0_184), .A1 (n_0_0_74), .A2 (n_0_0_183), .B1 (n_0_0_90), .B2 (n_0_0_171));
AOI22_X1 i_0_0_256 (.ZN (n_0_0_183), .A1 (n_0_0_182), .A2 (hfn_ipo_n64), .B1 (n_0_0_155), .B2 (hfn_ipo_n82));
OAI22_X1 i_0_0_255 (.ZN (n_0_0_182), .A1 (n_0_0_136), .A2 (hfn_ipo_n61), .B1 (n_0_0_181), .B2 (hfn_ipo_n79));
OAI22_X1 i_0_0_254 (.ZN (n_0_0_181), .A1 (n_0_0_140), .A2 (n_0_0_179), .B1 (n_0_0_86), .B2 (n_0_0_180));
INV_X1 i_0_0_253 (.ZN (n_0_0_180), .A (\extended_M[12] ));
INV_X1 i_0_0_252 (.ZN (n_0_0_179), .A (\extended_M[4] ));
AOI22_X1 i_0_0_251 (.ZN (n_0_0_178), .A1 (hfn_ipo_n66), .A2 (n_0_0_177), .B1 (n_0_0_94), .B2 (n_0_0_166));
OAI22_X1 i_0_0_250 (.ZN (n_0_0_177), .A1 (n_0_0_176), .A2 (hfn_ipo_n82), .B1 (n_0_0_160), .B2 (hfn_ipo_n64));
OAI22_X1 i_0_0_249 (.ZN (n_0_0_176), .A1 (n_0_0_131), .A2 (hfn_ipo_n61), .B1 (n_0_0_175), .B2 (hfn_ipo_n79));
OAI22_X1 i_0_0_248 (.ZN (n_0_0_175), .A1 (n_0_0_140), .A2 (n_0_0_173), .B1 (n_0_0_86), .B2 (n_0_0_174));
INV_X1 i_0_0_247 (.ZN (n_0_0_174), .A (\extended_M_mul_neg_one[12] ));
INV_X1 i_0_0_246 (.ZN (n_0_0_173), .A (\extended_M_mul_neg_one[4] ));
NAND2_X1 i_0_0_245 (.ZN (\partialProd[11] ), .A1 (n_0_0_167), .A2 (n_0_0_172));
AOI22_X1 i_0_0_244 (.ZN (n_0_0_172), .A1 (hfn_ipo_n66), .A2 (n_0_0_171), .B1 (n_0_0_90), .B2 (n_0_0_161));
OAI22_X1 i_0_0_243 (.ZN (n_0_0_171), .A1 (n_0_0_144), .A2 (hfn_ipo_n64), .B1 (n_0_0_170), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_0_242 (.ZN (n_0_0_170), .A1 (n_0_0_169), .A2 (hfn_ipo_n61), .B1 (n_0_0_17), .B2 (\extended_M_mul_neg_one[7] ));
OAI22_X1 i_0_0_241 (.ZN (n_0_0_169), .A1 (n_0_0_140), .A2 (n_0_0_96), .B1 (n_0_0_86), .B2 (n_0_0_168));
INV_X1 i_0_0_240 (.ZN (n_0_0_168), .A (\extended_M_mul_neg_one[11] ));
AOI22_X1 i_0_0_239 (.ZN (n_0_0_167), .A1 (n_0_0_74), .A2 (n_0_0_166), .B1 (n_0_0_94), .B2 (n_0_0_156));
OAI22_X1 i_0_0_238 (.ZN (n_0_0_166), .A1 (n_0_0_150), .A2 (hfn_ipo_n64), .B1 (n_0_0_165), .B2 (hfn_ipo_n82));
AOI22_X1 i_0_0_237 (.ZN (n_0_0_165), .A1 (n_0_0_164), .A2 (hfn_ipo_n61), .B1 (n_0_0_17), .B2 (\extended_M[7] ));
OAI22_X1 i_0_0_236 (.ZN (n_0_0_164), .A1 (n_0_0_140), .A2 (n_0_0_101), .B1 (n_0_0_86), .B2 (n_0_0_163));
INV_X1 i_0_0_235 (.ZN (n_0_0_163), .A (\extended_M[11] ));
NAND2_X1 i_0_0_234 (.ZN (\partialProd[10] ), .A1 (n_0_0_157), .A2 (n_0_0_162));
AOI22_X1 i_0_0_233 (.ZN (n_0_0_162), .A1 (hfn_ipo_n66), .A2 (n_0_0_161), .B1 (n_0_0_90), .B2 (n_0_0_145));
AOI22_X1 i_0_0_232 (.ZN (n_0_0_161), .A1 (n_0_0_132), .A2 (hfn_ipo_n82), .B1 (n_0_0_160), .B2 (hfn_ipo_n64));
AOI22_X1 i_0_0_231 (.ZN (n_0_0_160), .A1 (n_0_0_159), .A2 (hfn_ipo_n61), .B1 (\extended_M_mul_neg_one[6] ), .B2 (n_0_0_17));
OAI22_X1 i_0_0_230 (.ZN (n_0_0_159), .A1 (n_0_0_140), .A2 (n_0_0_114), .B1 (n_0_0_86), .B2 (n_0_0_158));
INV_X1 i_0_0_229 (.ZN (n_0_0_158), .A (\extended_M_mul_neg_one[10] ));
AOI22_X1 i_0_0_228 (.ZN (n_0_0_157), .A1 (n_0_0_74), .A2 (n_0_0_156), .B1 (n_0_0_94), .B2 (n_0_0_151));
OAI22_X1 i_0_0_227 (.ZN (n_0_0_156), .A1 (hfn_ipo_n82), .A2 (n_0_0_155), .B1 (n_0_0_137), .B2 (hfn_ipo_n64));
AOI22_X1 i_0_0_226 (.ZN (n_0_0_155), .A1 (n_0_0_154), .A2 (hfn_ipo_n61), .B1 (n_0_0_17), .B2 (\extended_M[6] ));
OAI22_X1 i_0_0_225 (.ZN (n_0_0_154), .A1 (n_0_0_140), .A2 (n_0_0_107), .B1 (n_0_0_86), .B2 (n_0_0_153));
INV_X1 i_0_0_224 (.ZN (n_0_0_153), .A (\extended_M[10] ));
NAND2_X1 i_0_0_223 (.ZN (\partialProd[9] ), .A1 (n_0_0_146), .A2 (n_0_0_152));
AOI22_X1 i_0_0_222 (.ZN (n_0_0_152), .A1 (n_0_0_74), .A2 (n_0_0_151), .B1 (n_0_0_90), .B2 (n_0_0_133));
OAI22_X1 i_0_0_221 (.ZN (n_0_0_151), .A1 (n_0_0_150), .A2 (hfn_ipo_n82), .B1 (hfn_ipo_n64), .B2 (n_0_0_122));
AOI22_X1 i_0_0_220 (.ZN (n_0_0_150), .A1 (n_0_0_149), .A2 (hfn_ipo_n61), .B1 (n_0_0_17), .B2 (\extended_M[5] ));
OAI22_X1 i_0_0_219 (.ZN (n_0_0_149), .A1 (n_0_0_140), .A2 (n_0_0_147), .B1 (n_0_0_86), .B2 (n_0_0_148));
INV_X1 i_0_0_218 (.ZN (n_0_0_148), .A (\extended_M[9] ));
INV_X1 i_0_0_217 (.ZN (n_0_0_147), .A (\extended_M[1] ));
AOI22_X1 i_0_0_216 (.ZN (n_0_0_146), .A1 (hfn_ipo_n66), .A2 (n_0_0_145), .B1 (n_0_0_94), .B2 (n_0_0_138));
OAI22_X1 i_0_0_215 (.ZN (n_0_0_145), .A1 (n_0_0_144), .A2 (hfn_ipo_n82), .B1 (n_0_0_100), .B2 (n_0_0_125));
AOI22_X1 i_0_0_214 (.ZN (n_0_0_144), .A1 (n_0_0_143), .A2 (hfn_ipo_n61), .B1 (n_0_0_17), .B2 (\extended_M_mul_neg_one[5] ));
OAI22_X1 i_0_0_213 (.ZN (n_0_0_143), .A1 (n_0_0_140), .A2 (n_0_0_141), .B1 (n_0_0_86), .B2 (n_0_0_142));
INV_X1 i_0_0_212 (.ZN (n_0_0_142), .A (\extended_M_mul_neg_one[9] ));
INV_X1 i_0_0_211 (.ZN (n_0_0_141), .A (\extended_M_mul_neg_one[1] ));
INV_X1 i_0_0_210 (.ZN (n_0_0_140), .A (n_0_0_128));
NAND2_X1 i_0_0_209 (.ZN (\partialProd[8] ), .A1 (n_0_0_134), .A2 (n_0_0_139));
AOI22_X1 i_0_0_208 (.ZN (n_0_0_139), .A1 (n_0_0_74), .A2 (n_0_0_138), .B1 (n_0_0_90), .B2 (n_0_0_126));
OAI22_X1 i_0_0_207 (.ZN (n_0_0_138), .A1 (n_0_0_137), .A2 (hfn_ipo_n82), .B1 (hfn_ipo_n64), .B2 (n_0_0_110));
AOI22_X1 i_0_0_206 (.ZN (n_0_0_137), .A1 (n_0_0_136), .A2 (hfn_ipo_n61), .B1 (\extended_M[4] ), .B2 (n_0_0_17));
OAI21_X1 i_0_0_205 (.ZN (n_0_0_136), .A (n_0_0_129), .B1 (n_0_0_135), .B2 (n_0_0_86));
INV_X1 i_0_0_204 (.ZN (n_0_0_135), .A (\extended_M[8] ));
AOI22_X1 i_0_0_203 (.ZN (n_0_0_134), .A1 (hfn_ipo_n66), .A2 (n_0_0_133), .B1 (n_0_0_94), .B2 (n_0_0_123));
OAI22_X1 i_0_0_202 (.ZN (n_0_0_133), .A1 (n_0_0_132), .A2 (hfn_ipo_n82), .B1 (n_0_0_117), .B2 (hfn_ipo_n64));
AOI22_X1 i_0_0_201 (.ZN (n_0_0_132), .A1 (n_0_0_131), .A2 (hfn_ipo_n61), .B1 (\extended_M_mul_neg_one[4] ), .B2 (n_0_0_17));
OAI21_X1 i_0_0_200 (.ZN (n_0_0_131), .A (n_0_0_129), .B1 (n_0_0_130), .B2 (n_0_0_86));
INV_X1 i_0_0_199 (.ZN (n_0_0_130), .A (\extended_M_mul_neg_one[8] ));
NAND2_X1 i_0_0_198 (.ZN (n_0_0_129), .A1 (n_0_0_128), .A2 (\extended_M[0] ));
NOR2_X2 i_0_0_197 (.ZN (n_0_0_128), .A1 (n_0_0_8), .A2 (drc_ipo_n83));
NAND2_X1 i_0_0_196 (.ZN (\partialProd[7] ), .A1 (n_0_0_124), .A2 (n_0_0_127));
AOI22_X1 i_0_0_195 (.ZN (n_0_0_127), .A1 (hfn_ipo_n66), .A2 (n_0_0_126), .B1 (n_0_0_90), .B2 (n_0_0_118));
OAI33_X1 i_0_0_194 (.ZN (n_0_0_126), .A1 (n_0_0_97), .A2 (hfn_ipo_n64), .A3 (n_0_0_86)
    , .B1 (n_0_0_86), .B2 (n_0_0_125), .B3 (hfn_ipo_n82));
AOI22_X1 i_0_0_193 (.ZN (n_0_0_125), .A1 (hfn_ipo_n61), .A2 (\extended_M_mul_neg_one[7] )
    , .B1 (\extended_M_mul_neg_one[3] ), .B2 (hfn_ipo_n79));
AOI22_X1 i_0_0_192 (.ZN (n_0_0_124), .A1 (n_0_0_74), .A2 (n_0_0_123), .B1 (n_0_0_94), .B2 (n_0_0_111));
OAI22_X1 i_0_0_191 (.ZN (n_0_0_123), .A1 (n_0_0_102), .A2 (n_0_0_100), .B1 (n_0_0_122), .B2 (hfn_ipo_n82));
NAND2_X1 i_0_0_190 (.ZN (n_0_0_122), .A1 (n_0_0_85), .A2 (n_0_0_121));
OAI22_X1 i_0_0_189 (.ZN (n_0_0_121), .A1 (n_0_0_101), .A2 (hfn_ipo_n61), .B1 (n_0_0_120), .B2 (hfn_ipo_n79));
INV_X1 i_0_0_188 (.ZN (n_0_0_120), .A (\extended_M[7] ));
NAND2_X1 i_0_0_187 (.ZN (\partialProd[6] ), .A1 (n_0_0_112), .A2 (n_0_0_119));
AOI22_X1 i_0_0_186 (.ZN (n_0_0_119), .A1 (hfn_ipo_n66), .A2 (n_0_0_118), .B1 (n_0_0_94), .B2 (n_0_0_103));
OAI22_X1 i_0_0_185 (.ZN (n_0_0_118), .A1 (n_0_0_100), .A2 (n_0_0_113), .B1 (n_0_0_117), .B2 (hfn_ipo_n82));
NAND2_X1 i_0_0_184 (.ZN (n_0_0_117), .A1 (n_0_0_85), .A2 (n_0_0_116));
OAI22_X1 i_0_0_183 (.ZN (n_0_0_116), .A1 (n_0_0_114), .A2 (hfn_ipo_n60), .B1 (n_0_0_115), .B2 (hfn_ipo_n79));
INV_X1 i_0_0_182 (.ZN (n_0_0_115), .A (\extended_M_mul_neg_one[6] ));
INV_X1 i_0_0_181 (.ZN (n_0_0_114), .A (\extended_M_mul_neg_one[2] ));
AOI22_X1 i_0_0_180 (.ZN (n_0_0_113), .A1 (hfn_ipo_n61), .A2 (\extended_M_mul_neg_one[4] )
    , .B1 (\extended_M[0] ), .B2 (hfn_ipo_n79));
AOI22_X1 i_0_0_179 (.ZN (n_0_0_112), .A1 (n_0_0_74), .A2 (n_0_0_111), .B1 (n_0_0_90), .B2 (n_0_0_98));
AOI21_X1 i_0_0_178 (.ZN (n_0_0_111), .A (n_0_0_106), .B1 (hfn_ipo_n64), .B2 (n_0_0_110));
NAND2_X1 i_0_0_177 (.ZN (n_0_0_110), .A1 (n_0_0_85), .A2 (n_0_0_109));
OAI22_X1 i_0_0_176 (.ZN (n_0_0_109), .A1 (n_0_0_107), .A2 (hfn_ipo_n61), .B1 (n_0_0_108), .B2 (hfn_ipo_n79));
INV_X1 i_0_0_175 (.ZN (n_0_0_108), .A (\extended_M[6] ));
INV_X1 i_0_0_174 (.ZN (n_0_0_107), .A (\extended_M[2] ));
AOI221_X1 i_0_0_173 (.ZN (n_0_0_106), .A (hfn_ipo_n64), .B1 (n_0_0_17), .B2 (\extended_M[0] )
    , .C1 (\extended_M[4] ), .C2 (n_0_0_105));
INV_X1 i_0_0_172 (.ZN (n_0_0_105), .A (n_0_0_57));
NAND2_X1 i_0_0_171 (.ZN (\partialProd[5] ), .A1 (n_0_0_99), .A2 (n_0_0_104));
AOI22_X1 i_0_0_170 (.ZN (n_0_0_104), .A1 (n_0_0_74), .A2 (n_0_0_103), .B1 (n_0_0_94), .B2 (n_0_0_93));
OAI33_X1 i_0_0_169 (.ZN (n_0_0_103), .A1 (n_0_0_100), .A2 (n_0_0_101), .A3 (hfn_ipo_n79)
    , .B1 (n_0_0_86), .B2 (n_0_0_102), .B3 (hfn_ipo_n82));
AOI22_X1 i_0_0_168 (.ZN (n_0_0_102), .A1 (hfn_ipo_n61), .A2 (\extended_M[5] ), .B1 (\extended_M[1] ), .B2 (hfn_ipo_n79));
INV_X1 i_0_0_167 (.ZN (n_0_0_101), .A (\extended_M[3] ));
NAND2_X1 i_0_0_166 (.ZN (n_0_0_100), .A1 (n_0_0_85), .A2 (hfn_ipo_n82));
AOI22_X1 i_0_0_165 (.ZN (n_0_0_99), .A1 (hfn_ipo_n66), .A2 (n_0_0_98), .B1 (n_0_0_90), .B2 (n_0_0_89));
OAI33_X1 i_0_0_164 (.ZN (n_0_0_98), .A1 (n_0_0_96), .A2 (hfn_ipo_n64), .A3 (n_0_0_57)
    , .B1 (n_0_0_86), .B2 (n_0_0_97), .B3 (hfn_ipo_n82));
AOI22_X1 i_0_0_163 (.ZN (n_0_0_97), .A1 (hfn_ipo_n61), .A2 (\extended_M_mul_neg_one[5] )
    , .B1 (\extended_M_mul_neg_one[1] ), .B2 (hfn_ipo_n79));
INV_X1 i_0_0_162 (.ZN (n_0_0_96), .A (\extended_M_mul_neg_one[3] ));
NAND2_X1 i_0_0_161 (.ZN (\partialProd[4] ), .A1 (n_0_0_91), .A2 (n_0_0_95));
AOI22_X1 i_0_0_160 (.ZN (n_0_0_95), .A1 (n_0_0_74), .A2 (n_0_0_93), .B1 (n_0_0_94), .B2 (n_0_0_83));
INV_X1 i_0_0_159 (.ZN (n_0_0_94), .A (n_0_0_70));
AOI21_X1 i_0_0_158 (.ZN (n_0_0_93), .A (n_0_0_86), .B1 (n_0_0_92), .B2 (n_0_0_88));
OAI221_X1 i_0_0_157 (.ZN (n_0_0_92), .A (hfn_ipo_n61), .B1 (\extended_M[4] ), .B2 (hfn_ipo_n81)
    , .C1 (\extended_M[2] ), .C2 (hfn_ipo_n63));
AOI22_X1 i_0_0_156 (.ZN (n_0_0_91), .A1 (hfn_ipo_n66), .A2 (n_0_0_89), .B1 (n_0_0_90), .B2 (n_0_0_81));
INV_X1 i_0_0_155 (.ZN (n_0_0_90), .A (n_0_0_69));
AOI21_X1 i_0_0_154 (.ZN (n_0_0_89), .A (n_0_0_86), .B1 (n_0_0_87), .B2 (n_0_0_88));
NAND3_X1 i_0_0_153 (.ZN (n_0_0_88), .A1 (hfn_ipo_n63), .A2 (\extended_M[0] ), .A3 (hfn_ipo_n79));
OAI221_X1 i_0_0_152 (.ZN (n_0_0_87), .A (hfn_ipo_n60), .B1 (\extended_M_mul_neg_one[4] )
    , .B2 (hfn_ipo_n81), .C1 (\extended_M_mul_neg_one[2] ), .C2 (hfn_ipo_n63));
INV_X1 i_0_0_151 (.ZN (n_0_0_86), .A (n_0_0_85));
NOR2_X1 i_0_0_150 (.ZN (n_0_0_85), .A1 (n_0_0_14), .A2 (drc_ipo_n83));
OAI221_X1 i_0_0_149 (.ZN (\partialProd[3] ), .A (n_0_0_84), .B1 (n_0_0_70), .B2 (n_0_0_78)
    , .C1 (n_0_0_69), .C2 (n_0_0_77));
AOI22_X1 i_0_0_148 (.ZN (n_0_0_84), .A1 (hfn_ipo_n66), .A2 (n_0_0_81), .B1 (n_0_0_74), .B2 (n_0_0_83));
NOR2_X1 i_0_0_147 (.ZN (n_0_0_83), .A1 (n_0_0_57), .A2 (n_0_0_82));
AOI22_X1 i_0_0_146 (.ZN (n_0_0_82), .A1 (hfn_ipo_n63), .A2 (\extended_M[3] ), .B1 (\extended_M[1] ), .B2 (hfn_ipo_n81));
NOR2_X1 i_0_0_145 (.ZN (n_0_0_81), .A1 (n_0_0_57), .A2 (n_0_0_80));
AOI22_X1 i_0_0_144 (.ZN (n_0_0_80), .A1 (hfn_ipo_n63), .A2 (\extended_M_mul_neg_one[3] )
    , .B1 (\extended_M_mul_neg_one[1] ), .B2 (hfn_ipo_n81));
OAI222_X1 i_0_0_143 (.ZN (\partialProd[2] ), .A1 (n_0_0_67), .A2 (n_0_0_77), .B1 (n_0_0_73)
    , .B2 (n_0_0_78), .C1 (n_0_0_69), .C2 (n_0_0_79));
NAND2_X1 i_0_0_142 (.ZN (n_0_0_79), .A1 (n_0_0_58), .A2 (\extended_M_mul_neg_one[1] ));
AOI21_X1 i_0_0_141 (.ZN (n_0_0_78), .A (n_0_0_76), .B1 (\extended_M[2] ), .B2 (n_0_0_58));
AOI21_X1 i_0_0_140 (.ZN (n_0_0_77), .A (n_0_0_76), .B1 (\extended_M_mul_neg_one[2] ), .B2 (n_0_0_58));
NOR3_X1 i_0_0_139 (.ZN (n_0_0_76), .A1 (n_0_0_57), .A2 (n_0_0_56), .A3 (hfn_ipo_n64));
AOI21_X1 i_0_0_138 (.ZN (\partialProd[1] ), .A (n_0_0_59), .B1 (n_0_0_72), .B2 (n_0_0_75));
NAND2_X1 i_0_0_137 (.ZN (n_0_0_75), .A1 (n_0_0_74), .A2 (\extended_M[1] ));
INV_X1 i_0_0_136 (.ZN (n_0_0_74), .A (n_0_0_73));
NAND2_X1 i_0_0_135 (.ZN (n_0_0_73), .A1 (n_0_0_60), .A2 (n_0_0_65));
AOI22_X1 i_0_0_134 (.ZN (n_0_0_72), .A1 (hfn_ipo_n66), .A2 (\extended_M_mul_neg_one[1] )
    , .B1 (n_0_0_71), .B2 (\extended_M[0] ));
NAND2_X1 i_0_0_133 (.ZN (n_0_0_71), .A1 (n_0_0_69), .A2 (n_0_0_70));
NAND3_X1 i_0_0_132 (.ZN (n_0_0_70), .A1 (n_0_0_65), .A2 (n_0_0_37), .A3 (n_0_0_54));
NAND3_X1 i_0_0_131 (.ZN (n_0_0_69), .A1 (n_0_0_36), .A2 (n_0_0_66), .A3 (n_0_0_53));
INV_X1 i_0_0_130 (.ZN (n_0_0_68), .A (n_0_0_67));
NAND2_X1 i_0_0_129 (.ZN (n_0_0_67), .A1 (n_0_0_60), .A2 (n_0_0_66));
INV_X1 i_0_0_128 (.ZN (n_0_0_66), .A (n_0_0_65));
AOI22_X1 i_0_0_127 (.ZN (n_0_0_65), .A1 (n_0_0_62), .A2 (n_0_0_64), .B1 (n_0_0_44), .B2 (hfn_ipo_n62));
AOI21_X1 i_0_0_126 (.ZN (n_0_0_64), .A (hfn_ipo_n62), .B1 (n_0_0_63), .B2 (n_0_0_29));
AOI22_X1 i_0_0_125 (.ZN (n_0_0_63), .A1 (\Q[32] ), .A2 (n_0_0_9), .B1 (n_0_0_10), .B2 (\Q[24] ));
AOI221_X1 i_0_0_124 (.ZN (n_0_0_62), .A (n_0_0_61), .B1 (n_0_0_33), .B2 (n_0_0_46)
    , .C1 (n_0_0_20), .C2 (n_0_0_50));
AOI221_X1 i_0_0_123 (.ZN (n_0_0_61), .A (n_0_0_16), .B1 (n_0_0_9), .B2 (\Q[16] ), .C1 (\Q[8] ), .C2 (n_0_0_10));
INV_X1 i_0_0_122 (.ZN (n_0_0_60), .A (n_0_0_55));
NOR3_X1 i_0_0_121 (.ZN (\partialProd[0] ), .A1 (n_0_0_55), .A2 (n_0_0_56), .A3 (n_0_0_59));
INV_X1 i_0_0_120 (.ZN (n_0_0_59), .A (n_0_0_58));
NOR2_X1 i_0_0_119 (.ZN (n_0_0_58), .A1 (n_0_0_57), .A2 (hfn_ipo_n82));
NAND2_X1 i_0_0_118 (.ZN (n_0_0_57), .A1 (n_0_0_20), .A2 (n_0_0_10));
INV_X1 i_0_0_117 (.ZN (n_0_0_56), .A (\extended_M[0] ));
OAI22_X1 i_0_0_116 (.ZN (n_0_0_55), .A1 (n_0_0_37), .A2 (n_0_0_54), .B1 (n_0_0_36), .B2 (n_0_0_53));
INV_X1 i_0_0_115 (.ZN (n_0_0_54), .A (n_0_0_53));
OAI22_X1 i_0_0_114 (.ZN (n_0_0_53), .A1 (n_0_0_44), .A2 (hfn_ipo_n62), .B1 (n_0_0_49), .B2 (n_0_0_52));
OAI22_X1 i_0_0_113 (.ZN (n_0_0_52), .A1 (n_0_0_50), .A2 (n_0_0_16), .B1 (n_0_0_51), .B2 (n_0_0_24));
AOI22_X1 i_0_0_112 (.ZN (n_0_0_51), .A1 (n_0_0_9), .A2 (\Q[24] ), .B1 (n_0_0_10), .B2 (\Q[16] ));
AOI22_X1 i_0_0_111 (.ZN (n_0_0_50), .A1 (n_0_0_9), .A2 (\Q[12] ), .B1 (n_0_0_10), .B2 (\Q[4] ));
OAI221_X1 i_0_0_110 (.ZN (n_0_0_49), .A (hfn_ipo_n62), .B1 (n_0_0_46), .B2 (n_0_0_12)
    , .C1 (n_0_0_48), .C2 (n_0_0_21));
AOI22_X1 i_0_0_109 (.ZN (n_0_0_48), .A1 (n_0_0_9), .A2 (\Q[8] ), .B1 (n_0_0_47), .B2 (\Q[32] ));
NOR2_X1 i_0_0_108 (.ZN (n_0_0_47), .A1 (n_0_0_7), .A2 (hfn_ipo_n75));
AOI22_X1 i_0_0_107 (.ZN (n_0_0_46), .A1 (n_0_0_9), .A2 (\Q[28] ), .B1 (n_0_0_10), .B2 (\Q[20] ));
INV_X1 i_0_0_106 (.ZN (n_0_0_45), .A (hfn_ipo_n81));
OAI211_X1 i_0_0_105 (.ZN (n_0_0_44), .A (n_0_0_41), .B (n_0_0_42), .C1 (n_0_0_24), .C2 (n_0_0_43));
AOI22_X1 i_0_0_104 (.ZN (n_0_0_43), .A1 (n_0_0_9), .A2 (\Q[26] ), .B1 (n_0_0_10), .B2 (\Q[18] ));
AOI22_X1 i_0_0_103 (.ZN (n_0_0_42), .A1 (\Q[6] ), .A2 (n_0_0_17), .B1 (n_0_0_18), .B2 (\Q[14] ));
INV_X1 i_0_0_102 (.ZN (n_0_0_41), .A (n_0_0_40));
OAI22_X1 i_0_0_101 (.ZN (n_0_0_40), .A1 (n_0_0_38), .A2 (n_0_0_12), .B1 (n_0_0_39), .B2 (n_0_0_21));
AOI22_X1 i_0_0_100 (.ZN (n_0_0_39), .A1 (n_0_0_9), .A2 (\Q[10] ), .B1 (n_0_0_10), .B2 (\Q[2] ));
AOI22_X1 i_0_0_99 (.ZN (n_0_0_38), .A1 (n_0_0_9), .A2 (\Q[30] ), .B1 (n_0_0_10), .B2 (\Q[22] ));
INV_X1 i_0_0_98 (.ZN (n_0_0_37), .A (n_0_0_36));
AOI22_X1 i_0_0_97 (.ZN (n_0_0_36), .A1 (n_0_0_26), .A2 (hfn_ipo_n80), .B1 (n_0_0_31), .B2 (n_0_0_35));
AOI22_X1 i_0_0_96 (.ZN (n_0_0_35), .A1 (n_0_0_32), .A2 (n_0_0_33), .B1 (n_0_0_34), .B2 (n_0_0_20));
AOI22_X1 i_0_0_95 (.ZN (n_0_0_34), .A1 (\Q[9] ), .A2 (n_0_0_9), .B1 (n_0_0_10), .B2 (\Q[1] ));
INV_X1 i_0_0_94 (.ZN (n_0_0_33), .A (n_0_0_24));
AOI22_X1 i_0_0_93 (.ZN (n_0_0_32), .A1 (\Q[25] ), .A2 (n_0_0_9), .B1 (n_0_0_10), .B2 (\Q[17] ));
AOI221_X1 i_0_0_92 (.ZN (n_0_0_31), .A (hfn_ipo_n80), .B1 (n_0_0_27), .B2 (n_0_0_28)
    , .C1 (n_0_0_29), .C2 (n_0_0_30));
AOI22_X1 i_0_0_91 (.ZN (n_0_0_30), .A1 (n_0_0_9), .A2 (\Q[29] ), .B1 (n_0_0_10), .B2 (\Q[21] ));
INV_X1 i_0_0_90 (.ZN (n_0_0_29), .A (n_0_0_12));
INV_X1 i_0_0_89 (.ZN (n_0_0_28), .A (n_0_0_16));
AOI22_X1 i_0_0_88 (.ZN (n_0_0_27), .A1 (\Q[13] ), .A2 (n_0_0_9), .B1 (n_0_0_10), .B2 (\Q[5] ));
OAI221_X1 i_0_0_87 (.ZN (n_0_0_26), .A (n_0_0_19), .B1 (n_0_0_21), .B2 (n_0_0_22)
    , .C1 (n_0_0_24), .C2 (n_0_0_25));
AOI22_X1 i_0_0_86 (.ZN (n_0_0_25), .A1 (n_0_0_9), .A2 (\Q[27] ), .B1 (n_0_0_10), .B2 (\Q[19] ));
NAND2_X1 i_0_0_85 (.ZN (n_0_0_24), .A1 (hfn_ipo_n59), .A2 (drc_ipo_n83));
INV_X1 i_0_0_84 (.ZN (n_0_0_23), .A (hfn_ipo_n78));
AOI22_X1 i_0_0_83 (.ZN (n_0_0_22), .A1 (n_0_0_9), .A2 (\Q[11] ), .B1 (n_0_0_10), .B2 (\Q[3] ));
INV_X1 i_0_0_82 (.ZN (n_0_0_21), .A (n_0_0_20));
NOR2_X1 i_0_0_81 (.ZN (n_0_0_20), .A1 (drc_ipo_n83), .A2 (hfn_ipo_n77));
AOI221_X1 i_0_0_80 (.ZN (n_0_0_19), .A (n_0_0_13), .B1 (\Q[7] ), .B2 (n_0_0_17), .C1 (\Q[15] ), .C2 (n_0_0_18));
NOR2_X1 i_0_0_79 (.ZN (n_0_0_18), .A1 (n_0_0_8), .A2 (n_0_0_16));
NOR2_X2 i_0_0_78 (.ZN (n_0_0_17), .A1 (n_0_0_14), .A2 (n_0_0_16));
NAND2_X1 i_0_0_77 (.ZN (n_0_0_16), .A1 (n_0_0_15), .A2 (hfn_ipo_n77));
INV_X2 i_0_0_76 (.ZN (n_0_0_15), .A (drc_ipo_n83));
INV_X1 i_0_0_75 (.ZN (n_0_0_14), .A (n_0_0_10));
NOR2_X1 i_0_0_74 (.ZN (n_0_0_13), .A1 (n_0_0_11), .A2 (n_0_0_12));
NAND2_X1 i_0_0_73 (.ZN (n_0_0_12), .A1 (drc_ipo_n83), .A2 (hfn_ipo_n77));
AOI22_X1 i_0_0_72 (.ZN (n_0_0_11), .A1 (n_0_0_9), .A2 (\Q[31] ), .B1 (n_0_0_10), .B2 (\Q[23] ));
NOR2_X4 i_0_0_71 (.ZN (n_0_0_10), .A1 (hfn_ipo_n75), .A2 (drc_ipo_n84));
INV_X1 i_0_0_70 (.ZN (n_0_0_9), .A (n_0_0_8));
NAND2_X1 i_0_0_69 (.ZN (n_0_0_8), .A1 (n_0_0_7), .A2 (hfn_ipo_n75));
INV_X2 i_0_0_68 (.ZN (n_0_0_7), .A (drc_ipo_n84));
AND2_X1 i_0_0_67 (.ZN (n_0_159), .A1 (n_0_0_6), .A2 (n_0_95));
AND2_X1 i_0_0_66 (.ZN (n_0_158), .A1 (n_0_0_6), .A2 (n_0_94));
AND2_X1 i_0_0_65 (.ZN (n_0_157), .A1 (n_0_0_6), .A2 (n_0_93));
AND2_X1 i_0_0_64 (.ZN (n_0_156), .A1 (n_0_0_6), .A2 (n_0_92));
AND2_X1 i_0_0_63 (.ZN (n_0_155), .A1 (n_0_0_6), .A2 (n_0_91));
AND2_X1 i_0_0_62 (.ZN (n_0_154), .A1 (n_0_0_6), .A2 (n_0_90));
AND2_X1 i_0_0_61 (.ZN (n_0_153), .A1 (n_0_0_6), .A2 (n_0_89));
AND2_X1 i_0_0_60 (.ZN (n_0_152), .A1 (n_0_0_6), .A2 (n_0_88));
AND2_X1 i_0_0_59 (.ZN (n_0_151), .A1 (n_0_0_6), .A2 (n_0_87));
AND2_X1 i_0_0_58 (.ZN (n_0_150), .A1 (n_0_0_6), .A2 (n_0_86));
AND2_X1 i_0_0_57 (.ZN (n_0_149), .A1 (n_0_0_6), .A2 (n_0_85));
AND2_X1 i_0_0_56 (.ZN (n_0_148), .A1 (n_0_0_6), .A2 (n_0_84));
AND2_X1 i_0_0_55 (.ZN (n_0_147), .A1 (n_0_0_6), .A2 (n_0_83));
AND2_X1 i_0_0_54 (.ZN (n_0_146), .A1 (n_0_0_6), .A2 (n_0_82));
AND2_X1 i_0_0_53 (.ZN (n_0_145), .A1 (n_0_0_6), .A2 (n_0_81));
AND2_X1 i_0_0_52 (.ZN (n_0_144), .A1 (n_0_0_6), .A2 (n_0_80));
AND2_X1 i_0_0_51 (.ZN (n_0_143), .A1 (n_0_0_6), .A2 (n_0_79));
AND2_X1 i_0_0_50 (.ZN (n_0_142), .A1 (n_0_0_6), .A2 (n_0_78));
AND2_X1 i_0_0_49 (.ZN (n_0_141), .A1 (n_0_0_6), .A2 (n_0_77));
AND2_X1 i_0_0_48 (.ZN (n_0_140), .A1 (n_0_0_6), .A2 (n_0_76));
AND2_X1 i_0_0_47 (.ZN (n_0_139), .A1 (n_0_0_6), .A2 (n_0_75));
AND2_X1 i_0_0_46 (.ZN (n_0_138), .A1 (n_0_0_6), .A2 (n_0_74));
AND2_X1 i_0_0_45 (.ZN (n_0_137), .A1 (n_0_0_6), .A2 (n_0_73));
AND2_X1 i_0_0_44 (.ZN (n_0_136), .A1 (n_0_0_6), .A2 (n_0_72));
AND2_X1 i_0_0_43 (.ZN (n_0_135), .A1 (hfn_ipo_n57), .A2 (n_0_71));
AND2_X1 i_0_0_42 (.ZN (n_0_134), .A1 (hfn_ipo_n57), .A2 (n_0_70));
AND2_X1 i_0_0_41 (.ZN (n_0_133), .A1 (hfn_ipo_n57), .A2 (n_0_69));
AND2_X1 i_0_0_40 (.ZN (n_0_132), .A1 (hfn_ipo_n57), .A2 (n_0_68));
AND2_X1 i_0_0_39 (.ZN (n_0_131), .A1 (hfn_ipo_n57), .A2 (n_0_67));
AND2_X1 i_0_0_38 (.ZN (n_0_130), .A1 (hfn_ipo_n57), .A2 (n_0_66));
AND2_X1 i_0_0_37 (.ZN (n_0_129), .A1 (hfn_ipo_n57), .A2 (n_0_65));
AND2_X1 i_0_0_36 (.ZN (n_0_128), .A1 (hfn_ipo_n57), .A2 (n_0_64));
AND2_X1 i_0_0_35 (.ZN (n_0_127), .A1 (hfn_ipo_n57), .A2 (n_0_63));
AND2_X1 i_0_0_34 (.ZN (n_0_126), .A1 (hfn_ipo_n57), .A2 (n_0_62));
AND2_X1 i_0_0_33 (.ZN (n_0_125), .A1 (hfn_ipo_n57), .A2 (n_0_61));
AND2_X1 i_0_0_32 (.ZN (n_0_124), .A1 (hfn_ipo_n57), .A2 (n_0_60));
AND2_X1 i_0_0_31 (.ZN (n_0_123), .A1 (hfn_ipo_n57), .A2 (n_0_59));
AND2_X1 i_0_0_30 (.ZN (n_0_122), .A1 (hfn_ipo_n57), .A2 (n_0_58));
AND2_X1 i_0_0_29 (.ZN (n_0_121), .A1 (hfn_ipo_n57), .A2 (n_0_57));
AND2_X1 i_0_0_28 (.ZN (n_0_120), .A1 (hfn_ipo_n57), .A2 (n_0_56));
AND2_X1 i_0_0_27 (.ZN (n_0_119), .A1 (hfn_ipo_n57), .A2 (n_0_55));
AND2_X1 i_0_0_26 (.ZN (n_0_118), .A1 (hfn_ipo_n57), .A2 (n_0_54));
AND2_X1 i_0_0_25 (.ZN (n_0_117), .A1 (hfn_ipo_n57), .A2 (n_0_53));
AND2_X1 i_0_0_24 (.ZN (n_0_116), .A1 (hfn_ipo_n57), .A2 (n_0_52));
AND2_X1 i_0_0_23 (.ZN (n_0_115), .A1 (hfn_ipo_n57), .A2 (n_0_51));
AND2_X1 i_0_0_22 (.ZN (n_0_114), .A1 (hfn_ipo_n57), .A2 (n_0_50));
AND2_X1 i_0_0_21 (.ZN (n_0_113), .A1 (hfn_ipo_n57), .A2 (n_0_49));
AND2_X1 i_0_0_20 (.ZN (n_0_112), .A1 (hfn_ipo_n57), .A2 (n_0_48));
AND2_X1 i_0_0_19 (.ZN (n_0_111), .A1 (hfn_ipo_n57), .A2 (n_0_47));
AND2_X1 i_0_0_18 (.ZN (n_0_110), .A1 (hfn_ipo_n57), .A2 (n_0_46));
AND2_X1 i_0_0_17 (.ZN (n_0_109), .A1 (hfn_ipo_n57), .A2 (n_0_45));
AND2_X1 i_0_0_16 (.ZN (n_0_108), .A1 (hfn_ipo_n57), .A2 (n_0_44));
AND2_X1 i_0_0_15 (.ZN (n_0_107), .A1 (hfn_ipo_n57), .A2 (n_0_43));
AND2_X1 i_0_0_14 (.ZN (n_0_106), .A1 (hfn_ipo_n57), .A2 (n_0_42));
AND2_X1 i_0_0_13 (.ZN (n_0_105), .A1 (hfn_ipo_n57), .A2 (n_0_41));
AND2_X1 i_0_0_12 (.ZN (n_0_104), .A1 (hfn_ipo_n57), .A2 (n_0_40));
AND2_X1 i_0_0_11 (.ZN (n_0_103), .A1 (hfn_ipo_n57), .A2 (n_0_39));
AND2_X1 i_0_0_10 (.ZN (n_0_102), .A1 (hfn_ipo_n57), .A2 (n_0_38));
AND2_X1 i_0_0_9 (.ZN (n_0_101), .A1 (hfn_ipo_n57), .A2 (n_0_37));
AND2_X1 i_0_0_8 (.ZN (n_0_100), .A1 (hfn_ipo_n57), .A2 (n_0_36));
AND2_X1 i_0_0_7 (.ZN (n_0_99), .A1 (hfn_ipo_n57), .A2 (n_0_35));
AND2_X1 i_0_0_6 (.ZN (n_0_98), .A1 (hfn_ipo_n57), .A2 (n_0_34));
AND2_X1 i_0_0_5 (.ZN (n_0_97), .A1 (hfn_ipo_n57), .A2 (n_0_33));
AND2_X1 i_0_0_4 (.ZN (n_0_96), .A1 (hfn_ipo_n57), .A2 (n_0_1));
INV_X1 i_0_0_3 (.ZN (n_0_0_6), .A (start));
HA_X1 i_0_0_2 (.CO (n_0_0_2), .S (n_0_0_5), .A (drc_ipo_n83), .B (n_0_0_1));
HA_X1 i_0_0_1 (.CO (n_0_0_1), .S (n_0_0_4), .A (hfn_ipo_n75), .B (n_0_0_0));
HA_X1 i_0_0_0 (.CO (n_0_0_0), .S (n_0_0_3), .A (hfn_ipo_n77), .B (hfn_ipo_n80));
datapath__0_19 i_0_14 (.p_0 ({n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, 
    n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, 
    n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, 
    n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, 
    n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, 
    n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, 
    n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_1}), .Acc ({\Acc[63] , \Acc[62] , 
    \Acc[61] , \Acc[60] , \Acc[59] , \Acc[58] , \Acc[57] , \Acc[56] , \Acc[55] , 
    \Acc[54] , \Acc[53] , \Acc[52] , \Acc[51] , \Acc[50] , \Acc[49] , \Acc[48] , 
    \Acc[47] , \Acc[46] , \Acc[45] , \Acc[44] , \Acc[43] , \Acc[42] , \Acc[41] , 
    \Acc[40] , \Acc[39] , \Acc[38] , \Acc[37] , \Acc[36] , \Acc[35] , \Acc[34] , 
    \Acc[33] , \Acc[32] , \Acc[31] , \Acc[30] , \Acc[29] , \Acc[28] , \Acc[27] , 
    \Acc[26] , \Acc[25] , \Acc[24] , \Acc[23] , \Acc[22] , \Acc[21] , \Acc[20] , 
    \Acc[19] , \Acc[18] , \Acc[17] , \Acc[16] , \Acc[15] , \Acc[14] , \Acc[13] , 
    \Acc[12] , \Acc[11] , \Acc[10] , \Acc[9] , \Acc[8] , \Acc[7] , \Acc[6] , \Acc[5] , 
    \Acc[4] , \Acc[3] , \Acc[2] , \Acc[1] , \Acc[0] }), .partialProd ({\partialProd[63] , 
    \partialProd[62] , \partialProd[61] , \partialProd[60] , \partialProd[59] , \partialProd[58] , 
    \partialProd[57] , \partialProd[56] , \partialProd[55] , \partialProd[54] , \partialProd[53] , 
    \partialProd[52] , \partialProd[51] , \partialProd[50] , \partialProd[49] , \partialProd[48] , 
    \partialProd[47] , \partialProd[46] , \partialProd[45] , \partialProd[44] , \partialProd[43] , 
    \partialProd[42] , \partialProd[41] , \partialProd[40] , \partialProd[39] , \partialProd[38] , 
    \partialProd[37] , \partialProd[36] , \partialProd[35] , \partialProd[34] , \partialProd[33] , 
    \partialProd[32] , \partialProd[31] , \partialProd[30] , \partialProd[29] , \partialProd[28] , 
    \partialProd[27] , \partialProd[26] , \partialProd[25] , \partialProd[24] , \partialProd[23] , 
    \partialProd[22] , \partialProd[21] , \partialProd[20] , \partialProd[19] , \partialProd[18] , 
    \partialProd[17] , \partialProd[16] , \partialProd[15] , \partialProd[14] , \partialProd[13] , 
    \partialProd[12] , \partialProd[11] , \partialProd[10] , \partialProd[9] , \partialProd[8] , 
    \partialProd[7] , \partialProd[6] , \partialProd[5] , \partialProd[4] , \partialProd[3] , 
    \partialProd[2] , \partialProd[1] , \partialProd[0] }));
datapath i_0_1 (.p_0 ({n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
    n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, 
    n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, 
    n_0_3, n_0_2, uc_0}), .A_reg ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }));
DFF_X1 \out_reg_reg[0]  (.Q (\out_reg[0] ), .CK (CTS_n214), .D (\Acc[0] ));
DFF_X1 \out_reg_reg[1]  (.Q (\out_reg[1] ), .CK (CTS_n214), .D (\Acc[1] ));
DFF_X1 \out_reg_reg[2]  (.Q (\out_reg[2] ), .CK (CTS_n214), .D (\Acc[2] ));
DFF_X1 \out_reg_reg[3]  (.Q (\out_reg[3] ), .CK (CTS_n214), .D (\Acc[3] ));
DFF_X1 \out_reg_reg[4]  (.Q (\out_reg[4] ), .CK (CTS_n214), .D (\Acc[4] ));
DFF_X1 \out_reg_reg[5]  (.Q (\out_reg[5] ), .CK (CTS_n214), .D (\Acc[5] ));
DFF_X1 \out_reg_reg[6]  (.Q (\out_reg[6] ), .CK (CTS_n214), .D (\Acc[6] ));
DFF_X1 \out_reg_reg[7]  (.Q (\out_reg[7] ), .CK (CTS_n214), .D (\Acc[7] ));
DFF_X1 \out_reg_reg[8]  (.Q (\out_reg[8] ), .CK (CTS_n214), .D (\Acc[8] ));
DFF_X1 \out_reg_reg[9]  (.Q (\out_reg[9] ), .CK (CTS_n214), .D (\Acc[9] ));
DFF_X1 \out_reg_reg[10]  (.Q (\out_reg[10] ), .CK (CTS_n214), .D (\Acc[10] ));
DFF_X1 \out_reg_reg[11]  (.Q (\out_reg[11] ), .CK (CTS_n214), .D (\Acc[11] ));
DFF_X1 \out_reg_reg[12]  (.Q (\out_reg[12] ), .CK (CTS_n214), .D (\Acc[12] ));
DFF_X1 \out_reg_reg[13]  (.Q (\out_reg[13] ), .CK (CTS_n214), .D (\Acc[13] ));
DFF_X1 \out_reg_reg[14]  (.Q (\out_reg[14] ), .CK (CTS_n214), .D (\Acc[14] ));
DFF_X1 \out_reg_reg[15]  (.Q (\out_reg[15] ), .CK (CTS_n214), .D (\Acc[15] ));
DFF_X1 \out_reg_reg[16]  (.Q (\out_reg[16] ), .CK (CTS_n214), .D (\Acc[16] ));
DFF_X1 \out_reg_reg[17]  (.Q (\out_reg[17] ), .CK (CTS_n214), .D (\Acc[17] ));
DFF_X1 \out_reg_reg[18]  (.Q (\out_reg[18] ), .CK (CTS_n214), .D (\Acc[18] ));
DFF_X1 \out_reg_reg[19]  (.Q (\out_reg[19] ), .CK (CTS_n214), .D (\Acc[19] ));
DFF_X1 \out_reg_reg[20]  (.Q (\out_reg[20] ), .CK (CTS_n214), .D (\Acc[20] ));
DFF_X1 \out_reg_reg[21]  (.Q (\out_reg[21] ), .CK (CTS_n214), .D (\Acc[21] ));
DFF_X1 \out_reg_reg[22]  (.Q (\out_reg[22] ), .CK (CTS_n214), .D (\Acc[22] ));
DFF_X1 \out_reg_reg[23]  (.Q (\out_reg[23] ), .CK (CTS_n214), .D (\Acc[23] ));
DFF_X1 \out_reg_reg[24]  (.Q (\out_reg[24] ), .CK (CTS_n214), .D (\Acc[24] ));
DFF_X1 \out_reg_reg[25]  (.Q (\out_reg[25] ), .CK (CTS_n214), .D (\Acc[25] ));
DFF_X1 \out_reg_reg[26]  (.Q (\out_reg[26] ), .CK (CTS_n214), .D (\Acc[26] ));
DFF_X1 \out_reg_reg[27]  (.Q (\out_reg[27] ), .CK (CTS_n214), .D (\Acc[27] ));
DFF_X1 \out_reg_reg[28]  (.Q (\out_reg[28] ), .CK (CTS_n214), .D (\Acc[28] ));
DFF_X1 \out_reg_reg[29]  (.Q (\out_reg[29] ), .CK (CTS_n214), .D (\Acc[29] ));
DFF_X1 \out_reg_reg[30]  (.Q (\out_reg[30] ), .CK (CTS_n214), .D (\Acc[30] ));
DFF_X1 \out_reg_reg[31]  (.Q (\out_reg[31] ), .CK (CTS_n214), .D (\Acc[31] ));
DFF_X1 \out_reg_reg[32]  (.Q (\out_reg[32] ), .CK (CTS_n214), .D (\Acc[32] ));
DFF_X1 \out_reg_reg[33]  (.Q (\out_reg[33] ), .CK (CTS_n214), .D (\Acc[33] ));
DFF_X1 \out_reg_reg[34]  (.Q (\out_reg[34] ), .CK (CTS_n214), .D (\Acc[34] ));
DFF_X1 \out_reg_reg[35]  (.Q (\out_reg[35] ), .CK (CTS_n214), .D (\Acc[35] ));
DFF_X1 \out_reg_reg[36]  (.Q (\out_reg[36] ), .CK (CTS_n214), .D (\Acc[36] ));
DFF_X1 \out_reg_reg[37]  (.Q (\out_reg[37] ), .CK (CTS_n214), .D (\Acc[37] ));
DFF_X1 \out_reg_reg[38]  (.Q (\out_reg[38] ), .CK (CTS_n214), .D (\Acc[38] ));
DFF_X1 \out_reg_reg[39]  (.Q (\out_reg[39] ), .CK (CTS_n214), .D (\Acc[39] ));
DFF_X1 \out_reg_reg[40]  (.Q (\out_reg[40] ), .CK (CTS_n214), .D (\Acc[40] ));
DFF_X1 \out_reg_reg[41]  (.Q (\out_reg[41] ), .CK (CTS_n214), .D (\Acc[41] ));
DFF_X1 \out_reg_reg[42]  (.Q (\out_reg[42] ), .CK (CTS_n214), .D (\Acc[42] ));
DFF_X1 \out_reg_reg[43]  (.Q (\out_reg[43] ), .CK (CTS_n214), .D (\Acc[43] ));
DFF_X1 \out_reg_reg[44]  (.Q (\out_reg[44] ), .CK (CTS_n214), .D (\Acc[44] ));
DFF_X1 \out_reg_reg[45]  (.Q (\out_reg[45] ), .CK (CTS_n214), .D (\Acc[45] ));
DFF_X1 \out_reg_reg[46]  (.Q (\out_reg[46] ), .CK (CTS_n214), .D (\Acc[46] ));
DFF_X1 \out_reg_reg[47]  (.Q (\out_reg[47] ), .CK (CTS_n214), .D (\Acc[47] ));
DFF_X1 \out_reg_reg[48]  (.Q (\out_reg[48] ), .CK (CTS_n214), .D (\Acc[48] ));
DFF_X1 \out_reg_reg[49]  (.Q (\out_reg[49] ), .CK (CTS_n214), .D (\Acc[49] ));
DFF_X1 \out_reg_reg[50]  (.Q (\out_reg[50] ), .CK (CTS_n214), .D (\Acc[50] ));
DFF_X1 \out_reg_reg[51]  (.Q (\out_reg[51] ), .CK (CTS_n214), .D (\Acc[51] ));
DFF_X1 \out_reg_reg[52]  (.Q (\out_reg[52] ), .CK (CTS_n214), .D (\Acc[52] ));
DFF_X1 \out_reg_reg[53]  (.Q (\out_reg[53] ), .CK (CTS_n214), .D (\Acc[53] ));
DFF_X1 \out_reg_reg[54]  (.Q (\out_reg[54] ), .CK (CTS_n214), .D (\Acc[54] ));
DFF_X1 \out_reg_reg[55]  (.Q (\out_reg[55] ), .CK (CTS_n214), .D (\Acc[55] ));
DFF_X1 \out_reg_reg[56]  (.Q (\out_reg[56] ), .CK (CTS_n214), .D (\Acc[56] ));
DFF_X1 \out_reg_reg[57]  (.Q (\out_reg[57] ), .CK (CTS_n214), .D (\Acc[57] ));
DFF_X1 \out_reg_reg[58]  (.Q (\out_reg[58] ), .CK (CTS_n214), .D (\Acc[58] ));
DFF_X1 \out_reg_reg[59]  (.Q (\out_reg[59] ), .CK (CTS_n214), .D (\Acc[59] ));
DFF_X1 \out_reg_reg[60]  (.Q (\out_reg[60] ), .CK (CTS_n214), .D (\Acc[60] ));
DFF_X1 \out_reg_reg[61]  (.Q (\out_reg[61] ), .CK (CTS_n214), .D (\Acc[61] ));
DFF_X1 \out_reg_reg[62]  (.Q (\out_reg[62] ), .CK (CTS_n214), .D (\Acc[62] ));
DFF_X1 \out_reg_reg[63]  (.Q (\out_reg[63] ), .CK (CTS_n214), .D (\Acc[63] ));
CLKGATETST_X8 clk_gate_out_reg_reg (.GCK (CTS_n215), .CK (CTS_n285), .E (n_0_166), .SE (VSS));
registerNbits__parameterized0 regOut (.out ({result[63], result[62], result[61], 
    result[60], result[59], result[58], result[57], result[56], result[55], result[54], 
    result[53], result[52], result[51], result[50], result[49], result[48], result[47], 
    result[46], result[45], result[44], result[43], result[42], result[41], result[40], 
    result[39], result[38], result[37], result[36], result[35], result[34], result[33], 
    result[32], result[31], result[30], result[29], result[28], result[27], result[26], 
    result[25], result[24], result[23], result[22], result[21], result[20], result[19], 
    result[18], result[17], result[16], result[15], result[14], result[13], result[12], 
    result[11], result[10], result[9], result[8], result[7], result[6], result[5], 
    result[4], result[3], result[2], result[1], result[0]}), .en (en), .inp ({\out_reg[63] , 
    \out_reg[62] , \out_reg[61] , \out_reg[60] , \out_reg[59] , \out_reg[58] , \out_reg[57] , 
    \out_reg[56] , \out_reg[55] , \out_reg[54] , \out_reg[53] , \out_reg[52] , \out_reg[51] , 
    \out_reg[50] , \out_reg[49] , \out_reg[48] , \out_reg[47] , \out_reg[46] , \out_reg[45] , 
    \out_reg[44] , \out_reg[43] , \out_reg[42] , \out_reg[41] , \out_reg[40] , \out_reg[39] , 
    \out_reg[38] , \out_reg[37] , \out_reg[36] , \out_reg[35] , \out_reg[34] , \out_reg[33] , 
    \out_reg[32] , \out_reg[31] , \out_reg[30] , \out_reg[29] , \out_reg[28] , \out_reg[27] , 
    \out_reg[26] , \out_reg[25] , \out_reg[24] , \out_reg[23] , \out_reg[22] , \out_reg[21] , 
    \out_reg[20] , \out_reg[19] , \out_reg[18] , \out_reg[17] , \out_reg[16] , \out_reg[15] , 
    \out_reg[14] , \out_reg[13] , \out_reg[12] , \out_reg[11] , \out_reg[10] , \out_reg[9] , 
    \out_reg[8] , \out_reg[7] , \out_reg[6] , \out_reg[5] , \out_reg[4] , \out_reg[3] , 
    \out_reg[2] , \out_reg[1] , \out_reg[0] }), .reset (reset), .clk_CTSPP_1 (CTS_n285));
registerNbits regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , \A_reg[27] , 
    \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , \A_reg[21] , 
    \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , \A_reg[15] , 
    \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , \A_reg[9] , 
    \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , 
    \A_reg[1] , \A_reg[0] }), .en (en), .inp ({inputA[31], inputA[30], inputA[29], 
    inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], inputA[22], 
    inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], inputA[15], 
    inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], inputA[8], 
    inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], inputA[1], 
    inputA[0]}), .reset (reset), .clk_CTSPP_1 (CTS_n285));
registerNbits__0_23 regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , 
    \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , 
    \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , 
    \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , 
    \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .en (en), .inp ({inputB[31], inputB[30], 
    inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], inputB[24], inputB[23], 
    inputB[22], inputB[21], inputB[20], inputB[19], inputB[18], inputB[17], inputB[16], 
    inputB[15], inputB[14], inputB[13], inputB[12], inputB[11], inputB[10], inputB[9], 
    inputB[8], inputB[7], inputB[6], inputB[5], inputB[4], inputB[3], inputB[2], 
    inputB[1], inputB[0]}), .reset (reset), .clk_CTSPP_1 (CTS_n285));
BUF_X2 hfn_ipo_c57 (.Z (hfn_ipo_n57), .A (n_0_0_6));
CLKBUF_X3 CTS_L3_c101 (.Z (CTS_n98), .A (CTS_n146));
CLKBUF_X3 CTS_L3_c102 (.Z (CTS_n99), .A (CTS_n146));
CLKBUF_X2 hfn_ipo_c75 (.Z (hfn_ipo_n75), .A (\i[3] ));
CLKBUF_X2 hfn_ipo_c76 (.Z (hfn_ipo_n76), .A (\i[3] ));
BUF_X4 hfn_ipo_c81 (.Z (hfn_ipo_n81), .A (\i[1] ));
BUF_X4 hfn_ipo_c82 (.Z (hfn_ipo_n82), .A (\i[1] ));
BUF_X4 drc_ipo_c83 (.Z (drc_ipo_n83), .A (\i[4] ));
BUF_X4 hfn_ipo_c59 (.Z (hfn_ipo_n59), .A (n_0_0_23));
BUF_X2 hfn_ipo_c60 (.Z (hfn_ipo_n60), .A (n_0_0_23));
CLKBUF_X2 hfn_ipo_c65 (.Z (hfn_ipo_n65), .A (n_0_0_68));
CLKBUF_X1 hfn_ipo_c66 (.Z (hfn_ipo_n66), .A (n_0_0_68));
BUF_X2 hfn_ipo_c61 (.Z (hfn_ipo_n61), .A (n_0_0_23));
BUF_X4 hfn_ipo_c62 (.Z (hfn_ipo_n62), .A (n_0_0_45));
BUF_X4 hfn_ipo_c63 (.Z (hfn_ipo_n63), .A (n_0_0_45));
BUF_X2 hfn_ipo_c64 (.Z (hfn_ipo_n64), .A (n_0_0_45));
CLKBUF_X1 CTS_L2_c2_c255 (.Z (CLOCK_n311), .A (CTS_n285));
CLKBUF_X1 hfn_ipo_c71 (.Z (hfn_ipo_n71), .A (n_0_0_94));
CLKBUF_X1 hfn_ipo_c69 (.Z (hfn_ipo_n69), .A (n_0_0_90));
CLKBUF_X3 CTS_L4_c189 (.Z (CTS_n188), .A (CTS_n187));
CLKBUF_X1 hfn_ipo_c73 (.Z (hfn_ipo_n73), .A (n_0_0_318));
BUF_X4 hfn_ipo_c77 (.Z (hfn_ipo_n77), .A (\i[2] ));
BUF_X2 hfn_ipo_c78 (.Z (hfn_ipo_n78), .A (\i[2] ));
BUF_X2 hfn_ipo_c79 (.Z (hfn_ipo_n79), .A (\i[2] ));
BUF_X4 hfn_ipo_c80 (.Z (hfn_ipo_n80), .A (\i[1] ));
BUF_X4 drc_ipo_c84 (.Z (drc_ipo_n84), .A (\i[5] ));
CLKBUF_X3 CTS_L4_c190 (.Z (CTS_n189), .A (CTS_n187));
CLKBUF_X1 hfn_ipo_c67 (.Z (hfn_ipo_n67), .A (n_0_0_74));
CLKBUF_X3 CTS_L4_c191 (.Z (CTS_n190), .A (CTS_n187));
CLKBUF_X1 CLOCK_slh__c266 (.Z (CLOCK_slh_n317), .A (start));
CLKBUF_X3 CTS_L3_c209 (.Z (CTS_n214), .A (CTS_n215));
CLKBUF_X3 CTS_L1_c1_c256 (.Z (CTS_n285), .A (clk));

endmodule //RadixBooth


