/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Jan  3 19:50:50 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1124999740 */

module datapath(p_0, p_1);
   output [31:0]p_0;
   input [31:0]p_1;

   XOR2_X1 i_0 (.A(p_1[1]), .B(p_1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(p_1[2]), .B1(p_1[1]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(p_1[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(p_1[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(p_1[6]), .B1(n_27), .B2(p_1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(p_1[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(p_1[9]), .B1(n_25), .B2(p_1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(p_1[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(p_1[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(p_1[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(p_1[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(p_1[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(p_1[16]), .B1(n_19), .B2(p_1[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(p_1[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(p_1[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(p_1[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(p_1[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(p_1[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(p_1[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(p_1[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(p_1[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(p_1[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(p_1[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(p_1[27]), .B1(n_9), .B2(p_1[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(p_1[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(p_1[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(p_1[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(p_1[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .A4(p_1[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(p_1[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(p_1[26]), .A3(p_1[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(p_1[23]), .A3(p_1[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(p_1[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(p_1[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .A4(p_1[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(p_1[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(p_1[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(p_1[15]), .A3(p_1[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(p_1[12]), .A3(p_1[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(p_1[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(p_1[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(p_1[8]), .A3(p_1[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(p_1[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(p_1[5]), .A3(p_1[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(p_1[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(p_1[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(p_1[2]), .A2(p_1[1]), .A3(p_1[0]), .ZN(n_29));
   INV_X1 i_61 (.A(p_1[11]), .ZN(n_30));
   INV_X1 i_62 (.A(p_1[14]), .ZN(n_31));
   INV_X1 i_63 (.A(p_1[21]), .ZN(n_32));
   INV_X1 i_64 (.A(p_1[25]), .ZN(n_33));
endmodule

module datapath__0_8(p_0, p_1);
   output [63:0]p_0;
   input [63:0]p_1;

   XOR2_X1 i_0 (.A(p_1[1]), .B(p_1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(p_1[2]), .B1(p_1[1]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_1[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(p_1[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(p_1[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(p_1[6]), .B1(n_27), .B2(p_1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_1[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(p_1[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(p_1[9]), .B1(n_25), .B2(p_1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_1[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(p_1[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(p_1[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(p_1[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(p_1[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(p_1[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(p_1[16]), .B1(n_19), .B2(p_1[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(p_1[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(p_1[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(p_1[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(p_1[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(p_1[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(p_1[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(p_1[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(p_1[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(p_1[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(p_1[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(p_1[27]), .B1(n_9), .B2(p_1[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(p_1[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(p_1[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(p_1[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(p_1[31]), .B(n_5), .ZN(p_0[31]));
   NOR2_X1 i_36 (.A1(p_1[31]), .A2(n_5), .ZN(p_0[63]));
   NOR4_X1 i_37 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .A4(p_1[30]), .ZN(n_5));
   NOR3_X1 i_38 (.A1(n_8), .A2(p_1[28]), .A3(p_1[29]), .ZN(n_6));
   NOR2_X1 i_39 (.A1(n_8), .A2(p_1[28]), .ZN(n_7));
   OR3_X1 i_40 (.A1(n_9), .A2(p_1[26]), .A3(p_1[27]), .ZN(n_8));
   NAND2_X1 i_41 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_42 (.A1(n_12), .A2(p_1[23]), .A3(p_1[24]), .ZN(n_10));
   NOR2_X1 i_43 (.A1(n_12), .A2(p_1[23]), .ZN(n_11));
   OR2_X1 i_44 (.A1(n_13), .A2(p_1[22]), .ZN(n_12));
   NAND2_X1 i_45 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_46 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .A4(p_1[20]), .ZN(n_14));
   NOR3_X1 i_47 (.A1(n_17), .A2(p_1[18]), .A3(p_1[19]), .ZN(n_15));
   NOR2_X1 i_48 (.A1(n_17), .A2(p_1[18]), .ZN(n_16));
   OR2_X1 i_49 (.A1(n_18), .A2(p_1[17]), .ZN(n_17));
   OR3_X1 i_50 (.A1(n_19), .A2(p_1[15]), .A3(p_1[16]), .ZN(n_18));
   NAND2_X1 i_51 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_52 (.A1(n_22), .A2(p_1[12]), .A3(p_1[13]), .ZN(n_20));
   NOR2_X1 i_53 (.A1(n_22), .A2(p_1[12]), .ZN(n_21));
   NAND2_X1 i_54 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_55 (.A1(n_24), .A2(p_1[10]), .ZN(n_23));
   OR3_X1 i_56 (.A1(n_25), .A2(p_1[8]), .A3(p_1[9]), .ZN(n_24));
   OR2_X1 i_57 (.A1(n_26), .A2(p_1[7]), .ZN(n_25));
   OR3_X1 i_58 (.A1(n_27), .A2(p_1[5]), .A3(p_1[6]), .ZN(n_26));
   OR2_X1 i_59 (.A1(n_28), .A2(p_1[4]), .ZN(n_27));
   OR2_X1 i_60 (.A1(n_29), .A2(p_1[3]), .ZN(n_28));
   OR3_X1 i_61 (.A1(p_1[2]), .A2(p_1[1]), .A3(p_1[0]), .ZN(n_29));
   INV_X1 i_62 (.A(p_1[11]), .ZN(n_30));
   INV_X1 i_63 (.A(p_1[14]), .ZN(n_31));
   INV_X1 i_64 (.A(p_1[21]), .ZN(n_32));
   INV_X1 i_65 (.A(p_1[25]), .ZN(n_33));
endmodule

module datapath__0_14(multiplicand, accumulator, p_0);
   input [63:0]multiplicand;
   input [63:0]accumulator;
   output [63:0]p_0;

   HA_X1 i_0 (.A(multiplicand[0]), .B(accumulator[0]), .CO(n_0), .S(p_0[0]));
   FA_X1 i_1 (.A(multiplicand[1]), .B(accumulator[1]), .CI(n_0), .CO(n_1), 
      .S(p_0[1]));
   FA_X1 i_2 (.A(multiplicand[2]), .B(accumulator[2]), .CI(n_1), .CO(n_2), 
      .S(p_0[2]));
   FA_X1 i_3 (.A(multiplicand[3]), .B(accumulator[3]), .CI(n_2), .CO(n_3), 
      .S(p_0[3]));
   FA_X1 i_4 (.A(multiplicand[4]), .B(accumulator[4]), .CI(n_3), .CO(n_4), 
      .S(p_0[4]));
   FA_X1 i_5 (.A(multiplicand[5]), .B(accumulator[5]), .CI(n_4), .CO(n_5), 
      .S(p_0[5]));
   FA_X1 i_6 (.A(multiplicand[6]), .B(accumulator[6]), .CI(n_5), .CO(n_6), 
      .S(p_0[6]));
   FA_X1 i_7 (.A(multiplicand[7]), .B(accumulator[7]), .CI(n_6), .CO(n_7), 
      .S(p_0[7]));
   FA_X1 i_8 (.A(multiplicand[8]), .B(accumulator[8]), .CI(n_7), .CO(n_8), 
      .S(p_0[8]));
   FA_X1 i_9 (.A(multiplicand[9]), .B(accumulator[9]), .CI(n_8), .CO(n_9), 
      .S(p_0[9]));
   FA_X1 i_10 (.A(multiplicand[10]), .B(accumulator[10]), .CI(n_9), .CO(n_10), 
      .S(p_0[10]));
   FA_X1 i_11 (.A(multiplicand[11]), .B(accumulator[11]), .CI(n_10), .CO(n_11), 
      .S(p_0[11]));
   FA_X1 i_12 (.A(multiplicand[12]), .B(accumulator[12]), .CI(n_11), .CO(n_12), 
      .S(p_0[12]));
   FA_X1 i_13 (.A(multiplicand[13]), .B(accumulator[13]), .CI(n_12), .CO(n_13), 
      .S(p_0[13]));
   FA_X1 i_14 (.A(multiplicand[14]), .B(accumulator[14]), .CI(n_13), .CO(n_14), 
      .S(p_0[14]));
   FA_X1 i_15 (.A(multiplicand[15]), .B(accumulator[15]), .CI(n_14), .CO(n_15), 
      .S(p_0[15]));
   FA_X1 i_16 (.A(multiplicand[16]), .B(accumulator[16]), .CI(n_15), .CO(n_16), 
      .S(p_0[16]));
   FA_X1 i_17 (.A(multiplicand[17]), .B(accumulator[17]), .CI(n_16), .CO(n_17), 
      .S(p_0[17]));
   FA_X1 i_18 (.A(multiplicand[18]), .B(accumulator[18]), .CI(n_17), .CO(n_18), 
      .S(p_0[18]));
   FA_X1 i_19 (.A(multiplicand[19]), .B(accumulator[19]), .CI(n_18), .CO(n_19), 
      .S(p_0[19]));
   FA_X1 i_20 (.A(multiplicand[20]), .B(accumulator[20]), .CI(n_19), .CO(n_20), 
      .S(p_0[20]));
   FA_X1 i_21 (.A(multiplicand[21]), .B(accumulator[21]), .CI(n_20), .CO(n_21), 
      .S(p_0[21]));
   FA_X1 i_22 (.A(multiplicand[22]), .B(accumulator[22]), .CI(n_21), .CO(n_22), 
      .S(p_0[22]));
   FA_X1 i_23 (.A(multiplicand[23]), .B(accumulator[23]), .CI(n_22), .CO(n_23), 
      .S(p_0[23]));
   FA_X1 i_24 (.A(multiplicand[24]), .B(accumulator[24]), .CI(n_23), .CO(n_24), 
      .S(p_0[24]));
   FA_X1 i_25 (.A(multiplicand[25]), .B(accumulator[25]), .CI(n_24), .CO(n_25), 
      .S(p_0[25]));
   FA_X1 i_26 (.A(multiplicand[26]), .B(accumulator[26]), .CI(n_25), .CO(n_26), 
      .S(p_0[26]));
   FA_X1 i_27 (.A(multiplicand[27]), .B(accumulator[27]), .CI(n_26), .CO(n_27), 
      .S(p_0[27]));
   FA_X1 i_28 (.A(multiplicand[28]), .B(accumulator[28]), .CI(n_27), .CO(n_28), 
      .S(p_0[28]));
   FA_X1 i_29 (.A(multiplicand[29]), .B(accumulator[29]), .CI(n_28), .CO(n_29), 
      .S(p_0[29]));
   FA_X1 i_30 (.A(multiplicand[30]), .B(accumulator[30]), .CI(n_29), .CO(n_30), 
      .S(p_0[30]));
   FA_X1 i_31 (.A(multiplicand[31]), .B(accumulator[31]), .CI(n_30), .CO(n_31), 
      .S(p_0[31]));
   FA_X1 i_32 (.A(multiplicand[32]), .B(accumulator[32]), .CI(n_31), .CO(n_32), 
      .S(p_0[32]));
   FA_X1 i_33 (.A(multiplicand[33]), .B(accumulator[33]), .CI(n_32), .CO(n_33), 
      .S(p_0[33]));
   FA_X1 i_34 (.A(multiplicand[34]), .B(accumulator[34]), .CI(n_33), .CO(n_34), 
      .S(p_0[34]));
   FA_X1 i_35 (.A(multiplicand[35]), .B(accumulator[35]), .CI(n_34), .CO(n_35), 
      .S(p_0[35]));
   FA_X1 i_36 (.A(multiplicand[36]), .B(accumulator[36]), .CI(n_35), .CO(n_36), 
      .S(p_0[36]));
   FA_X1 i_37 (.A(multiplicand[37]), .B(accumulator[37]), .CI(n_36), .CO(n_37), 
      .S(p_0[37]));
   FA_X1 i_38 (.A(multiplicand[38]), .B(accumulator[38]), .CI(n_37), .CO(n_38), 
      .S(p_0[38]));
   FA_X1 i_39 (.A(multiplicand[39]), .B(accumulator[39]), .CI(n_38), .CO(n_39), 
      .S(p_0[39]));
   FA_X1 i_40 (.A(multiplicand[40]), .B(accumulator[40]), .CI(n_39), .CO(n_40), 
      .S(p_0[40]));
   FA_X1 i_41 (.A(multiplicand[41]), .B(accumulator[41]), .CI(n_40), .CO(n_41), 
      .S(p_0[41]));
   FA_X1 i_42 (.A(multiplicand[42]), .B(accumulator[42]), .CI(n_41), .CO(n_42), 
      .S(p_0[42]));
   FA_X1 i_43 (.A(multiplicand[43]), .B(accumulator[43]), .CI(n_42), .CO(n_43), 
      .S(p_0[43]));
   FA_X1 i_44 (.A(multiplicand[44]), .B(accumulator[44]), .CI(n_43), .CO(n_44), 
      .S(p_0[44]));
   FA_X1 i_45 (.A(multiplicand[45]), .B(accumulator[45]), .CI(n_44), .CO(n_45), 
      .S(p_0[45]));
   FA_X1 i_46 (.A(multiplicand[46]), .B(accumulator[46]), .CI(n_45), .CO(n_46), 
      .S(p_0[46]));
   FA_X1 i_47 (.A(multiplicand[47]), .B(accumulator[47]), .CI(n_46), .CO(n_47), 
      .S(p_0[47]));
   FA_X1 i_48 (.A(multiplicand[48]), .B(accumulator[48]), .CI(n_47), .CO(n_48), 
      .S(p_0[48]));
   FA_X1 i_49 (.A(multiplicand[49]), .B(accumulator[49]), .CI(n_48), .CO(n_49), 
      .S(p_0[49]));
   FA_X1 i_50 (.A(multiplicand[50]), .B(accumulator[50]), .CI(n_49), .CO(n_50), 
      .S(p_0[50]));
   FA_X1 i_51 (.A(multiplicand[51]), .B(accumulator[51]), .CI(n_50), .CO(n_51), 
      .S(p_0[51]));
   FA_X1 i_52 (.A(multiplicand[52]), .B(accumulator[52]), .CI(n_51), .CO(n_52), 
      .S(p_0[52]));
   FA_X1 i_53 (.A(multiplicand[53]), .B(accumulator[53]), .CI(n_52), .CO(n_53), 
      .S(p_0[53]));
   FA_X1 i_54 (.A(multiplicand[54]), .B(accumulator[54]), .CI(n_53), .CO(n_54), 
      .S(p_0[54]));
   FA_X1 i_55 (.A(multiplicand[55]), .B(accumulator[55]), .CI(n_54), .CO(n_55), 
      .S(p_0[55]));
   FA_X1 i_56 (.A(multiplicand[56]), .B(accumulator[56]), .CI(n_55), .CO(n_56), 
      .S(p_0[56]));
   FA_X1 i_57 (.A(multiplicand[57]), .B(accumulator[57]), .CI(n_56), .CO(n_57), 
      .S(p_0[57]));
   FA_X1 i_58 (.A(multiplicand[58]), .B(accumulator[58]), .CI(n_57), .CO(n_58), 
      .S(p_0[58]));
   FA_X1 i_59 (.A(multiplicand[59]), .B(accumulator[59]), .CI(n_58), .CO(n_59), 
      .S(p_0[59]));
   FA_X1 i_60 (.A(multiplicand[60]), .B(accumulator[60]), .CI(n_59), .CO(n_60), 
      .S(p_0[60]));
   FA_X1 i_61 (.A(multiplicand[61]), .B(accumulator[61]), .CI(n_60), .CO(n_61), 
      .S(p_0[61]));
   FA_X1 i_62 (.A(multiplicand[62]), .B(accumulator[62]), .CI(n_61), .CO(n_62), 
      .S(p_0[62]));
   XNOR2_X1 i_63 (.A(multiplicand[63]), .B(accumulator[63]), .ZN(n_63));
   XNOR2_X1 i_64 (.A(n_63), .B(n_62), .ZN(p_0[63]));
endmodule

module sequential_multiplier(clk, rst, x, y, product);
   input clk;
   input rst;
   input [31:0]x;
   input [31:0]y;
   output [63:0]product;

   wire n_0_0;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_0_3;
   wire n_0_0_0;
   wire n_0_0_4;
   wire n_0_0_1;
   wire n_0_0_5;
   wire n_0_0_2;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_0_8;
   wire n_0_212;
   wire n_0_0_9;
   wire n_0_213;
   wire n_0_0_10;
   wire n_0_214;
   wire n_0_0_11;
   wire n_0_215;
   wire n_0_0_12;
   wire n_0_216;
   wire n_0_0_13;
   wire n_0_217;
   wire n_0_0_14;
   wire n_0_218;
   wire n_0_0_15;
   wire n_0_219;
   wire n_0_0_16;
   wire n_0_220;
   wire n_0_0_17;
   wire n_0_221;
   wire n_0_0_18;
   wire n_0_222;
   wire n_0_0_19;
   wire n_0_223;
   wire n_0_0_20;
   wire n_0_224;
   wire n_0_0_21;
   wire n_0_225;
   wire n_0_0_22;
   wire n_0_226;
   wire n_0_0_23;
   wire n_0_227;
   wire n_0_0_24;
   wire n_0_228;
   wire n_0_0_25;
   wire n_0_229;
   wire n_0_0_26;
   wire n_0_230;
   wire n_0_0_27;
   wire n_0_231;
   wire n_0_0_28;
   wire n_0_232;
   wire n_0_0_29;
   wire n_0_233;
   wire n_0_0_30;
   wire n_0_234;
   wire n_0_0_31;
   wire n_0_235;
   wire n_0_0_32;
   wire n_0_236;
   wire n_0_0_33;
   wire n_0_237;
   wire n_0_0_34;
   wire n_0_238;
   wire n_0_0_35;
   wire n_0_239;
   wire n_0_0_36;
   wire n_0_240;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_241;
   wire n_0_0_39;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_0_40;
   wire n_0_274;
   wire n_0_275;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_0_79;
   wire n_0_371;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_372;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire [31:0]multiplier;
   wire [5:0]ctr;
   wire n_0_373;

   CLKGATETST_X1 clk_gate_product_reg (.CK(clk), .E(n_0_371), .SE(1'b0), 
      .GCK(n_0_0));
   DFF_X1 \product_reg[63]  (.D(n_0_375), .CK(n_0_0), .Q(product[63]), .QN());
   DFF_X1 \product_reg[62]  (.D(n_0_376), .CK(n_0_0), .Q(product[62]), .QN());
   DFF_X1 \product_reg[61]  (.D(n_0_377), .CK(n_0_0), .Q(product[61]), .QN());
   DFF_X1 \product_reg[60]  (.D(n_0_378), .CK(n_0_0), .Q(product[60]), .QN());
   DFF_X1 \product_reg[59]  (.D(n_0_379), .CK(n_0_0), .Q(product[59]), .QN());
   DFF_X1 \product_reg[58]  (.D(n_0_380), .CK(n_0_0), .Q(product[58]), .QN());
   DFF_X1 \product_reg[57]  (.D(n_0_381), .CK(n_0_0), .Q(product[57]), .QN());
   DFF_X1 \product_reg[56]  (.D(n_0_382), .CK(n_0_0), .Q(product[56]), .QN());
   DFF_X1 \product_reg[55]  (.D(n_0_383), .CK(n_0_0), .Q(product[55]), .QN());
   DFF_X1 \product_reg[54]  (.D(n_0_384), .CK(n_0_0), .Q(product[54]), .QN());
   DFF_X1 \product_reg[53]  (.D(n_0_385), .CK(n_0_0), .Q(product[53]), .QN());
   DFF_X1 \product_reg[52]  (.D(n_0_386), .CK(n_0_0), .Q(product[52]), .QN());
   DFF_X1 \product_reg[51]  (.D(n_0_387), .CK(n_0_0), .Q(product[51]), .QN());
   DFF_X1 \product_reg[50]  (.D(n_0_388), .CK(n_0_0), .Q(product[50]), .QN());
   DFF_X1 \product_reg[49]  (.D(n_0_389), .CK(n_0_0), .Q(product[49]), .QN());
   DFF_X1 \product_reg[48]  (.D(n_0_390), .CK(n_0_0), .Q(product[48]), .QN());
   DFF_X1 \product_reg[47]  (.D(n_0_391), .CK(n_0_0), .Q(product[47]), .QN());
   DFF_X1 \product_reg[46]  (.D(n_0_392), .CK(n_0_0), .Q(product[46]), .QN());
   DFF_X1 \product_reg[45]  (.D(n_0_393), .CK(n_0_0), .Q(product[45]), .QN());
   DFF_X1 \product_reg[44]  (.D(n_0_394), .CK(n_0_0), .Q(product[44]), .QN());
   DFF_X1 \product_reg[43]  (.D(n_0_395), .CK(n_0_0), .Q(product[43]), .QN());
   DFF_X1 \product_reg[42]  (.D(n_0_396), .CK(n_0_0), .Q(product[42]), .QN());
   DFF_X1 \product_reg[41]  (.D(n_0_397), .CK(n_0_0), .Q(product[41]), .QN());
   DFF_X1 \product_reg[40]  (.D(n_0_398), .CK(n_0_0), .Q(product[40]), .QN());
   DFF_X1 \product_reg[39]  (.D(n_0_399), .CK(n_0_0), .Q(product[39]), .QN());
   DFF_X1 \product_reg[38]  (.D(n_0_400), .CK(n_0_0), .Q(product[38]), .QN());
   DFF_X1 \product_reg[37]  (.D(n_0_401), .CK(n_0_0), .Q(product[37]), .QN());
   DFF_X1 \product_reg[36]  (.D(n_0_402), .CK(n_0_0), .Q(product[36]), .QN());
   DFF_X1 \product_reg[35]  (.D(n_0_403), .CK(n_0_0), .Q(product[35]), .QN());
   DFF_X1 \product_reg[34]  (.D(n_0_404), .CK(n_0_0), .Q(product[34]), .QN());
   DFF_X1 \product_reg[33]  (.D(n_0_405), .CK(n_0_0), .Q(product[33]), .QN());
   DFF_X1 \product_reg[32]  (.D(n_0_406), .CK(n_0_0), .Q(product[32]), .QN());
   DFF_X1 \product_reg[31]  (.D(n_0_407), .CK(n_0_0), .Q(product[31]), .QN());
   DFF_X1 \product_reg[30]  (.D(n_0_408), .CK(n_0_0), .Q(product[30]), .QN());
   DFF_X1 \product_reg[29]  (.D(n_0_409), .CK(n_0_0), .Q(product[29]), .QN());
   DFF_X1 \product_reg[28]  (.D(n_0_410), .CK(n_0_0), .Q(product[28]), .QN());
   DFF_X1 \product_reg[27]  (.D(n_0_411), .CK(n_0_0), .Q(product[27]), .QN());
   DFF_X1 \product_reg[26]  (.D(n_0_412), .CK(n_0_0), .Q(product[26]), .QN());
   DFF_X1 \product_reg[25]  (.D(n_0_413), .CK(n_0_0), .Q(product[25]), .QN());
   DFF_X1 \product_reg[24]  (.D(n_0_414), .CK(n_0_0), .Q(product[24]), .QN());
   DFF_X1 \product_reg[23]  (.D(n_0_415), .CK(n_0_0), .Q(product[23]), .QN());
   DFF_X1 \product_reg[22]  (.D(n_0_416), .CK(n_0_0), .Q(product[22]), .QN());
   DFF_X1 \product_reg[21]  (.D(n_0_417), .CK(n_0_0), .Q(product[21]), .QN());
   DFF_X1 \product_reg[20]  (.D(n_0_418), .CK(n_0_0), .Q(product[20]), .QN());
   DFF_X1 \product_reg[19]  (.D(n_0_419), .CK(n_0_0), .Q(product[19]), .QN());
   DFF_X1 \product_reg[18]  (.D(n_0_420), .CK(n_0_0), .Q(product[18]), .QN());
   DFF_X1 \product_reg[17]  (.D(n_0_421), .CK(n_0_0), .Q(product[17]), .QN());
   DFF_X1 \product_reg[16]  (.D(n_0_422), .CK(n_0_0), .Q(product[16]), .QN());
   DFF_X1 \product_reg[15]  (.D(n_0_423), .CK(n_0_0), .Q(product[15]), .QN());
   DFF_X1 \product_reg[14]  (.D(n_0_424), .CK(n_0_0), .Q(product[14]), .QN());
   DFF_X1 \product_reg[13]  (.D(n_0_425), .CK(n_0_0), .Q(product[13]), .QN());
   DFF_X1 \product_reg[12]  (.D(n_0_426), .CK(n_0_0), .Q(product[12]), .QN());
   DFF_X1 \product_reg[11]  (.D(n_0_427), .CK(n_0_0), .Q(product[11]), .QN());
   DFF_X1 \product_reg[10]  (.D(n_0_1), .CK(n_0_0), .Q(product[10]), .QN());
   DFF_X1 \product_reg[9]  (.D(n_0_2), .CK(n_0_0), .Q(product[9]), .QN());
   DFF_X1 \product_reg[8]  (.D(n_0_3), .CK(n_0_0), .Q(product[8]), .QN());
   DFF_X1 \product_reg[7]  (.D(n_0_4), .CK(n_0_0), .Q(product[7]), .QN());
   DFF_X1 \product_reg[6]  (.D(n_0_5), .CK(n_0_0), .Q(product[6]), .QN());
   DFF_X1 \product_reg[5]  (.D(n_0_6), .CK(n_0_0), .Q(product[5]), .QN());
   DFF_X1 \product_reg[4]  (.D(n_0_7), .CK(n_0_0), .Q(product[4]), .QN());
   DFF_X1 \product_reg[3]  (.D(n_0_8), .CK(n_0_0), .Q(product[3]), .QN());
   DFF_X1 \product_reg[2]  (.D(n_0_9), .CK(n_0_0), .Q(product[2]), .QN());
   DFF_X1 \product_reg[1]  (.D(n_0_10), .CK(n_0_0), .Q(product[1]), .QN());
   DFF_X1 \product_reg[0]  (.D(n_0_11), .CK(n_0_0), .Q(product[0]), .QN());
   datapath i_0_3 (.p_0({n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, 
      n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, 
      n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, 
      n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, uc_0}), .p_1({n_0_370, 
      n_0_369, n_0_368, n_0_367, n_0_366, n_0_365, n_0_364, n_0_363, n_0_362, 
      n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, n_0_356, n_0_355, n_0_354, 
      n_0_353, n_0_352, n_0_351, n_0_350, n_0_349, n_0_348, n_0_347, n_0_346, 
      n_0_345, n_0_344, n_0_343, n_0_342, n_0_341, n_0_340, n_0_339}));
   datapath__0_8 i_0_10 (.p_0({n_0_75, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, 
      uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, 
      uc_29, uc_30, uc_31, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, 
      n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, 
      n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, 
      n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, uc_32}), .p_1({
      uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, 
      uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, 
      uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, 
      uc_63, uc_64, n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, 
      n_0_332, n_0_331, n_0_330, n_0_329, n_0_328, n_0_327, n_0_326, n_0_325, 
      n_0_324, n_0_323, n_0_322, n_0_321, n_0_320, n_0_319, n_0_318, n_0_317, 
      n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, n_0_311, n_0_310, n_0_309, 
      n_0_308, n_0_307}));
   datapath__0_14 i_0_16 (.multiplicand({n_0_372, n_0_428, n_0_429, n_0_430, 
      n_0_431, n_0_432, n_0_433, n_0_434, n_0_435, n_0_436, n_0_437, n_0_438, 
      n_0_439, n_0_440, n_0_441, n_0_442, n_0_443, n_0_444, n_0_445, n_0_446, 
      n_0_447, n_0_448, n_0_449, n_0_450, n_0_451, n_0_452, n_0_453, n_0_454, 
      n_0_455, n_0_456, n_0_457, n_0_458, n_0_459, n_0_460, n_0_461, n_0_462, 
      n_0_463, n_0_464, n_0_465, n_0_466, n_0_467, n_0_468, n_0_469, n_0_470, 
      n_0_471, n_0_472, n_0_473, n_0_474, n_0_475, n_0_476, n_0_477, n_0_478, 
      n_0_479, n_0_480, n_0_481, n_0_482, n_0_483, n_0_484, n_0_485, n_0_486, 
      n_0_487, n_0_488, n_0_489, n_0_490}), .accumulator({n_0_375, n_0_376, 
      n_0_377, n_0_378, n_0_379, n_0_380, n_0_381, n_0_382, n_0_383, n_0_384, 
      n_0_385, n_0_386, n_0_387, n_0_388, n_0_389, n_0_390, n_0_391, n_0_392, 
      n_0_393, n_0_394, n_0_395, n_0_396, n_0_397, n_0_398, n_0_399, n_0_400, 
      n_0_401, n_0_402, n_0_403, n_0_404, n_0_405, n_0_406, n_0_407, n_0_408, 
      n_0_409, n_0_410, n_0_411, n_0_412, n_0_413, n_0_414, n_0_415, n_0_416, 
      n_0_417, n_0_418, n_0_419, n_0_420, n_0_421, n_0_422, n_0_423, n_0_424, 
      n_0_425, n_0_426, n_0_427, n_0_1, n_0_2, n_0_3, n_0_4, n_0_5, n_0_6, n_0_7, 
      n_0_8, n_0_9, n_0_10, n_0_11}), .p_0({n_0_139, n_0_138, n_0_137, n_0_136, 
      n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, 
      n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, 
      n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, 
      n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, 
      n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, 
      n_0_76}));
   HA_X1 i_0_0_0 (.A(ctr[1]), .B(ctr[0]), .CO(n_0_0_0), .S(n_0_0_3));
   HA_X1 i_0_0_1 (.A(ctr[2]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_4));
   HA_X1 i_0_0_2 (.A(ctr[3]), .B(n_0_0_1), .CO(n_0_0_2), .S(n_0_0_5));
   HA_X1 i_0_0_3 (.A(ctr[4]), .B(n_0_0_2), .CO(n_0_0_7), .S(n_0_0_6));
   AND2_X1 i_0_0_4 (.A1(n_0_0_119), .A2(n_0_76), .ZN(n_0_140));
   AND2_X1 i_0_0_5 (.A1(n_0_0_119), .A2(n_0_77), .ZN(n_0_141));
   AND2_X1 i_0_0_6 (.A1(n_0_0_119), .A2(n_0_78), .ZN(n_0_142));
   AND2_X1 i_0_0_7 (.A1(n_0_0_119), .A2(n_0_79), .ZN(n_0_143));
   AND2_X1 i_0_0_8 (.A1(n_0_0_119), .A2(n_0_80), .ZN(n_0_144));
   AND2_X1 i_0_0_9 (.A1(n_0_0_119), .A2(n_0_81), .ZN(n_0_145));
   AND2_X1 i_0_0_10 (.A1(n_0_0_119), .A2(n_0_82), .ZN(n_0_146));
   AND2_X1 i_0_0_11 (.A1(n_0_0_119), .A2(n_0_83), .ZN(n_0_147));
   AND2_X1 i_0_0_12 (.A1(n_0_0_119), .A2(n_0_84), .ZN(n_0_148));
   AND2_X1 i_0_0_13 (.A1(n_0_0_119), .A2(n_0_85), .ZN(n_0_149));
   AND2_X1 i_0_0_14 (.A1(n_0_0_119), .A2(n_0_86), .ZN(n_0_150));
   AND2_X1 i_0_0_15 (.A1(n_0_0_119), .A2(n_0_87), .ZN(n_0_151));
   AND2_X1 i_0_0_16 (.A1(n_0_0_119), .A2(n_0_88), .ZN(n_0_152));
   AND2_X1 i_0_0_17 (.A1(n_0_0_119), .A2(n_0_89), .ZN(n_0_153));
   AND2_X1 i_0_0_18 (.A1(n_0_0_119), .A2(n_0_90), .ZN(n_0_154));
   AND2_X1 i_0_0_19 (.A1(n_0_0_119), .A2(n_0_91), .ZN(n_0_155));
   AND2_X1 i_0_0_20 (.A1(n_0_0_119), .A2(n_0_92), .ZN(n_0_156));
   AND2_X1 i_0_0_21 (.A1(n_0_0_119), .A2(n_0_93), .ZN(n_0_157));
   AND2_X1 i_0_0_22 (.A1(n_0_0_119), .A2(n_0_94), .ZN(n_0_158));
   AND2_X1 i_0_0_23 (.A1(n_0_0_119), .A2(n_0_95), .ZN(n_0_159));
   AND2_X1 i_0_0_24 (.A1(n_0_0_119), .A2(n_0_96), .ZN(n_0_160));
   AND2_X1 i_0_0_25 (.A1(n_0_0_119), .A2(n_0_97), .ZN(n_0_161));
   AND2_X1 i_0_0_26 (.A1(n_0_0_119), .A2(n_0_98), .ZN(n_0_162));
   AND2_X1 i_0_0_27 (.A1(n_0_0_119), .A2(n_0_99), .ZN(n_0_163));
   AND2_X1 i_0_0_28 (.A1(n_0_0_119), .A2(n_0_100), .ZN(n_0_164));
   AND2_X1 i_0_0_29 (.A1(n_0_0_119), .A2(n_0_101), .ZN(n_0_165));
   AND2_X1 i_0_0_30 (.A1(n_0_0_119), .A2(n_0_102), .ZN(n_0_166));
   AND2_X1 i_0_0_31 (.A1(n_0_0_119), .A2(n_0_103), .ZN(n_0_167));
   AND2_X1 i_0_0_32 (.A1(n_0_0_119), .A2(n_0_104), .ZN(n_0_168));
   AND2_X1 i_0_0_33 (.A1(n_0_0_119), .A2(n_0_105), .ZN(n_0_169));
   AND2_X1 i_0_0_34 (.A1(n_0_0_119), .A2(n_0_106), .ZN(n_0_170));
   AND2_X1 i_0_0_35 (.A1(n_0_0_119), .A2(n_0_107), .ZN(n_0_171));
   AND2_X1 i_0_0_36 (.A1(n_0_0_119), .A2(n_0_108), .ZN(n_0_172));
   AND2_X1 i_0_0_37 (.A1(n_0_0_119), .A2(n_0_109), .ZN(n_0_173));
   AND2_X1 i_0_0_38 (.A1(n_0_0_119), .A2(n_0_110), .ZN(n_0_174));
   AND2_X1 i_0_0_39 (.A1(n_0_0_119), .A2(n_0_111), .ZN(n_0_175));
   AND2_X1 i_0_0_40 (.A1(n_0_0_119), .A2(n_0_112), .ZN(n_0_176));
   AND2_X1 i_0_0_41 (.A1(n_0_0_119), .A2(n_0_113), .ZN(n_0_177));
   AND2_X1 i_0_0_42 (.A1(n_0_0_119), .A2(n_0_114), .ZN(n_0_178));
   AND2_X1 i_0_0_43 (.A1(n_0_0_119), .A2(n_0_115), .ZN(n_0_179));
   AND2_X1 i_0_0_44 (.A1(n_0_0_119), .A2(n_0_116), .ZN(n_0_180));
   AND2_X1 i_0_0_45 (.A1(n_0_0_119), .A2(n_0_117), .ZN(n_0_181));
   AND2_X1 i_0_0_46 (.A1(n_0_0_119), .A2(n_0_118), .ZN(n_0_182));
   AND2_X1 i_0_0_47 (.A1(n_0_0_119), .A2(n_0_119), .ZN(n_0_183));
   AND2_X1 i_0_0_48 (.A1(n_0_0_119), .A2(n_0_120), .ZN(n_0_184));
   AND2_X1 i_0_0_49 (.A1(n_0_0_119), .A2(n_0_121), .ZN(n_0_185));
   AND2_X1 i_0_0_50 (.A1(n_0_0_119), .A2(n_0_122), .ZN(n_0_186));
   AND2_X1 i_0_0_51 (.A1(n_0_0_119), .A2(n_0_123), .ZN(n_0_187));
   AND2_X1 i_0_0_52 (.A1(n_0_0_119), .A2(n_0_124), .ZN(n_0_188));
   AND2_X1 i_0_0_53 (.A1(n_0_0_119), .A2(n_0_125), .ZN(n_0_189));
   AND2_X1 i_0_0_54 (.A1(n_0_0_119), .A2(n_0_126), .ZN(n_0_190));
   AND2_X1 i_0_0_55 (.A1(n_0_0_119), .A2(n_0_127), .ZN(n_0_191));
   AND2_X1 i_0_0_56 (.A1(n_0_0_119), .A2(n_0_128), .ZN(n_0_192));
   AND2_X1 i_0_0_57 (.A1(n_0_0_119), .A2(n_0_129), .ZN(n_0_193));
   AND2_X1 i_0_0_58 (.A1(n_0_0_119), .A2(n_0_130), .ZN(n_0_194));
   AND2_X1 i_0_0_59 (.A1(n_0_0_119), .A2(n_0_131), .ZN(n_0_195));
   AND2_X1 i_0_0_60 (.A1(n_0_0_119), .A2(n_0_132), .ZN(n_0_196));
   AND2_X1 i_0_0_61 (.A1(n_0_0_119), .A2(n_0_133), .ZN(n_0_197));
   AND2_X1 i_0_0_62 (.A1(n_0_0_119), .A2(n_0_134), .ZN(n_0_198));
   AND2_X1 i_0_0_63 (.A1(n_0_0_119), .A2(n_0_135), .ZN(n_0_199));
   AND2_X1 i_0_0_64 (.A1(n_0_0_119), .A2(n_0_136), .ZN(n_0_200));
   AND2_X1 i_0_0_65 (.A1(n_0_0_119), .A2(n_0_137), .ZN(n_0_201));
   AND2_X1 i_0_0_66 (.A1(n_0_0_119), .A2(n_0_138), .ZN(n_0_202));
   AND2_X1 i_0_0_67 (.A1(n_0_0_119), .A2(n_0_139), .ZN(n_0_203));
   NOR2_X1 i_0_0_68 (.A1(rst), .A2(ctr[0]), .ZN(n_0_204));
   AND2_X1 i_0_0_69 (.A1(n_0_0_119), .A2(n_0_0_3), .ZN(n_0_205));
   AND2_X1 i_0_0_70 (.A1(n_0_0_119), .A2(n_0_0_4), .ZN(n_0_206));
   AND2_X1 i_0_0_71 (.A1(n_0_0_119), .A2(n_0_0_5), .ZN(n_0_207));
   AND2_X1 i_0_0_72 (.A1(n_0_0_119), .A2(n_0_0_6), .ZN(n_0_208));
   AND2_X1 i_0_0_73 (.A1(n_0_0_119), .A2(n_0_0_7), .ZN(n_0_209));
   AND2_X1 i_0_0_74 (.A1(n_0_307), .A2(rst), .ZN(n_0_210));
   INV_X1 i_0_0_75 (.A(n_0_0_8), .ZN(n_0_211));
   AOI222_X1 i_0_0_76 (.A1(n_0_308), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_44), 
      .C1(n_0_0_80), .C2(n_0_490), .ZN(n_0_0_8));
   INV_X1 i_0_0_77 (.A(n_0_0_9), .ZN(n_0_212));
   AOI222_X1 i_0_0_78 (.A1(n_0_309), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_45), 
      .C1(n_0_0_80), .C2(n_0_489), .ZN(n_0_0_9));
   INV_X1 i_0_0_79 (.A(n_0_0_10), .ZN(n_0_213));
   AOI222_X1 i_0_0_80 (.A1(n_0_310), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_46), 
      .C1(n_0_0_80), .C2(n_0_488), .ZN(n_0_0_10));
   INV_X1 i_0_0_81 (.A(n_0_0_11), .ZN(n_0_214));
   AOI222_X1 i_0_0_82 (.A1(n_0_311), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_47), 
      .C1(n_0_0_80), .C2(n_0_487), .ZN(n_0_0_11));
   INV_X1 i_0_0_83 (.A(n_0_0_12), .ZN(n_0_215));
   AOI222_X1 i_0_0_84 (.A1(n_0_312), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_48), 
      .C1(n_0_0_80), .C2(n_0_486), .ZN(n_0_0_12));
   INV_X1 i_0_0_85 (.A(n_0_0_13), .ZN(n_0_216));
   AOI222_X1 i_0_0_86 (.A1(n_0_313), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_49), 
      .C1(n_0_0_80), .C2(n_0_485), .ZN(n_0_0_13));
   INV_X1 i_0_0_87 (.A(n_0_0_14), .ZN(n_0_217));
   AOI222_X1 i_0_0_88 (.A1(n_0_314), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_50), 
      .C1(n_0_0_80), .C2(n_0_484), .ZN(n_0_0_14));
   INV_X1 i_0_0_89 (.A(n_0_0_15), .ZN(n_0_218));
   AOI222_X1 i_0_0_90 (.A1(n_0_315), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_51), 
      .C1(n_0_0_80), .C2(n_0_483), .ZN(n_0_0_15));
   INV_X1 i_0_0_91 (.A(n_0_0_16), .ZN(n_0_219));
   AOI222_X1 i_0_0_92 (.A1(n_0_316), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_52), 
      .C1(n_0_0_80), .C2(n_0_482), .ZN(n_0_0_16));
   INV_X1 i_0_0_93 (.A(n_0_0_17), .ZN(n_0_220));
   AOI222_X1 i_0_0_94 (.A1(n_0_317), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_53), 
      .C1(n_0_0_80), .C2(n_0_481), .ZN(n_0_0_17));
   INV_X1 i_0_0_95 (.A(n_0_0_18), .ZN(n_0_221));
   AOI222_X1 i_0_0_96 (.A1(n_0_318), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_54), 
      .C1(n_0_0_80), .C2(n_0_480), .ZN(n_0_0_18));
   INV_X1 i_0_0_97 (.A(n_0_0_19), .ZN(n_0_222));
   AOI222_X1 i_0_0_98 (.A1(n_0_319), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_55), 
      .C1(n_0_0_80), .C2(n_0_479), .ZN(n_0_0_19));
   INV_X1 i_0_0_99 (.A(n_0_0_20), .ZN(n_0_223));
   AOI222_X1 i_0_0_100 (.A1(n_0_320), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_56), 
      .C1(n_0_0_80), .C2(n_0_478), .ZN(n_0_0_20));
   INV_X1 i_0_0_101 (.A(n_0_0_21), .ZN(n_0_224));
   AOI222_X1 i_0_0_102 (.A1(n_0_321), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_57), 
      .C1(n_0_0_80), .C2(n_0_477), .ZN(n_0_0_21));
   INV_X1 i_0_0_103 (.A(n_0_0_22), .ZN(n_0_225));
   AOI222_X1 i_0_0_104 (.A1(n_0_322), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_58), 
      .C1(n_0_0_80), .C2(n_0_476), .ZN(n_0_0_22));
   INV_X1 i_0_0_105 (.A(n_0_0_23), .ZN(n_0_226));
   AOI222_X1 i_0_0_106 (.A1(n_0_323), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_59), 
      .C1(n_0_0_80), .C2(n_0_475), .ZN(n_0_0_23));
   INV_X1 i_0_0_107 (.A(n_0_0_24), .ZN(n_0_227));
   AOI222_X1 i_0_0_108 (.A1(n_0_324), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_60), 
      .C1(n_0_0_80), .C2(n_0_474), .ZN(n_0_0_24));
   INV_X1 i_0_0_109 (.A(n_0_0_25), .ZN(n_0_228));
   AOI222_X1 i_0_0_110 (.A1(n_0_325), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_61), 
      .C1(n_0_0_80), .C2(n_0_473), .ZN(n_0_0_25));
   INV_X1 i_0_0_111 (.A(n_0_0_26), .ZN(n_0_229));
   AOI222_X1 i_0_0_112 (.A1(n_0_326), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_62), 
      .C1(n_0_0_80), .C2(n_0_472), .ZN(n_0_0_26));
   INV_X1 i_0_0_113 (.A(n_0_0_27), .ZN(n_0_230));
   AOI222_X1 i_0_0_114 (.A1(n_0_327), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_63), 
      .C1(n_0_0_80), .C2(n_0_471), .ZN(n_0_0_27));
   INV_X1 i_0_0_115 (.A(n_0_0_28), .ZN(n_0_231));
   AOI222_X1 i_0_0_116 (.A1(n_0_328), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_64), 
      .C1(n_0_0_80), .C2(n_0_470), .ZN(n_0_0_28));
   INV_X1 i_0_0_117 (.A(n_0_0_29), .ZN(n_0_232));
   AOI222_X1 i_0_0_118 (.A1(n_0_329), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_65), 
      .C1(n_0_0_80), .C2(n_0_469), .ZN(n_0_0_29));
   INV_X1 i_0_0_119 (.A(n_0_0_30), .ZN(n_0_233));
   AOI222_X1 i_0_0_120 (.A1(n_0_330), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_66), 
      .C1(n_0_0_80), .C2(n_0_468), .ZN(n_0_0_30));
   INV_X1 i_0_0_121 (.A(n_0_0_31), .ZN(n_0_234));
   AOI222_X1 i_0_0_122 (.A1(n_0_331), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_67), 
      .C1(n_0_0_80), .C2(n_0_467), .ZN(n_0_0_31));
   INV_X1 i_0_0_123 (.A(n_0_0_32), .ZN(n_0_235));
   AOI222_X1 i_0_0_124 (.A1(n_0_332), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_68), 
      .C1(n_0_0_80), .C2(n_0_466), .ZN(n_0_0_32));
   INV_X1 i_0_0_125 (.A(n_0_0_33), .ZN(n_0_236));
   AOI222_X1 i_0_0_126 (.A1(n_0_333), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_69), 
      .C1(n_0_0_80), .C2(n_0_465), .ZN(n_0_0_33));
   INV_X1 i_0_0_127 (.A(n_0_0_34), .ZN(n_0_237));
   AOI222_X1 i_0_0_128 (.A1(n_0_334), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_70), 
      .C1(n_0_0_80), .C2(n_0_464), .ZN(n_0_0_34));
   INV_X1 i_0_0_129 (.A(n_0_0_35), .ZN(n_0_238));
   AOI222_X1 i_0_0_130 (.A1(n_0_335), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_71), 
      .C1(n_0_0_80), .C2(n_0_463), .ZN(n_0_0_35));
   INV_X1 i_0_0_131 (.A(n_0_0_36), .ZN(n_0_239));
   AOI222_X1 i_0_0_132 (.A1(n_0_336), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_72), 
      .C1(n_0_0_80), .C2(n_0_462), .ZN(n_0_0_36));
   INV_X1 i_0_0_133 (.A(n_0_0_37), .ZN(n_0_240));
   AOI222_X1 i_0_0_134 (.A1(n_0_337), .A2(n_0_0_38), .B1(n_0_0_78), .B2(n_0_73), 
      .C1(n_0_0_80), .C2(n_0_461), .ZN(n_0_0_37));
   NOR2_X1 i_0_0_135 (.A1(n_0_370), .A2(n_0_0_119), .ZN(n_0_0_38));
   AOI21_X1 i_0_0_136 (.A(n_0_0_39), .B1(n_0_0_78), .B2(n_0_0_81), .ZN(n_0_241));
   AOI22_X1 i_0_0_137 (.A1(n_0_338), .A2(rst), .B1(n_0_460), .B2(n_0_0_80), 
      .ZN(n_0_0_39));
   OAI21_X1 i_0_0_138 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_82), .ZN(n_0_242));
   OAI21_X1 i_0_0_139 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_83), .ZN(n_0_243));
   OAI21_X1 i_0_0_140 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_84), .ZN(n_0_244));
   OAI21_X1 i_0_0_141 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_85), .ZN(n_0_245));
   OAI21_X1 i_0_0_142 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_86), .ZN(n_0_246));
   OAI21_X1 i_0_0_143 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_87), .ZN(n_0_247));
   OAI21_X1 i_0_0_144 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_88), .ZN(n_0_248));
   OAI21_X1 i_0_0_145 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_89), .ZN(n_0_249));
   OAI21_X1 i_0_0_146 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_90), .ZN(n_0_250));
   OAI21_X1 i_0_0_147 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_91), .ZN(n_0_251));
   OAI21_X1 i_0_0_148 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_92), .ZN(n_0_252));
   OAI21_X1 i_0_0_149 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_93), .ZN(n_0_253));
   OAI21_X1 i_0_0_150 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_94), .ZN(n_0_254));
   OAI21_X1 i_0_0_151 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_95), .ZN(n_0_255));
   OAI21_X1 i_0_0_152 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_96), .ZN(n_0_256));
   OAI21_X1 i_0_0_153 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_97), .ZN(n_0_257));
   OAI21_X1 i_0_0_154 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_98), .ZN(n_0_258));
   OAI21_X1 i_0_0_155 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_99), .ZN(n_0_259));
   OAI21_X1 i_0_0_156 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_100), .ZN(n_0_260));
   OAI21_X1 i_0_0_157 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_101), .ZN(n_0_261));
   OAI21_X1 i_0_0_158 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_102), .ZN(n_0_262));
   OAI21_X1 i_0_0_159 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_103), .ZN(n_0_263));
   OAI21_X1 i_0_0_160 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_104), .ZN(n_0_264));
   OAI21_X1 i_0_0_161 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_105), .ZN(n_0_265));
   OAI21_X1 i_0_0_162 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_106), .ZN(n_0_266));
   OAI21_X1 i_0_0_163 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_107), .ZN(n_0_267));
   OAI21_X1 i_0_0_164 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_108), .ZN(n_0_268));
   OAI21_X1 i_0_0_165 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_109), .ZN(n_0_269));
   OAI21_X1 i_0_0_166 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_110), .ZN(n_0_270));
   OAI21_X1 i_0_0_167 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_111), .ZN(n_0_271));
   OAI21_X1 i_0_0_168 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_112), .ZN(n_0_272));
   OAI21_X1 i_0_0_169 (.A(n_0_0_40), .B1(n_0_371), .B2(n_0_0_113), .ZN(n_0_273));
   OAI211_X1 i_0_0_170 (.A(n_0_338), .B(rst), .C1(n_0_75), .C2(n_0_0_79), 
      .ZN(n_0_0_40));
   NAND2_X1 i_0_0_171 (.A1(n_0_0_119), .A2(ctr[5]), .ZN(n_0_274));
   OAI21_X1 i_0_0_172 (.A(n_0_0_119), .B1(n_0_0_41), .B2(ctr[5]), .ZN(n_0_275));
   OAI21_X1 i_0_0_173 (.A(n_0_0_42), .B1(n_0_0_58), .B2(ctr[4]), .ZN(n_0_0_41));
   OAI221_X1 i_0_0_174 (.A(ctr[4]), .B1(n_0_0_50), .B2(n_0_0_43), .C1(n_0_0_51), 
      .C2(ctr[3]), .ZN(n_0_0_42));
   OAI221_X1 i_0_0_175 (.A(n_0_0_45), .B1(n_0_0_44), .B2(n_0_0_76), .C1(n_0_0_70), 
      .C2(multiplier[31]), .ZN(n_0_0_43));
   MUX2_X1 i_0_0_176 (.A(multiplier[24]), .B(multiplier[25]), .S(ctr[0]), 
      .Z(n_0_0_44));
   AOI22_X1 i_0_0_177 (.A1(n_0_0_49), .A2(n_0_0_48), .B1(n_0_0_47), .B2(n_0_0_46), 
      .ZN(n_0_0_45));
   AOI21_X1 i_0_0_178 (.A(n_0_0_75), .B1(multiplier[29]), .B2(ctr[0]), .ZN(
      n_0_0_46));
   NAND2_X1 i_0_0_179 (.A1(n_0_0_117), .A2(multiplier[28]), .ZN(n_0_0_47));
   AOI21_X1 i_0_0_180 (.A(n_0_0_74), .B1(multiplier[26]), .B2(n_0_0_117), 
      .ZN(n_0_0_48));
   NAND2_X1 i_0_0_181 (.A1(ctr[0]), .A2(multiplier[27]), .ZN(n_0_0_49));
   OAI21_X1 i_0_0_182 (.A(ctr[3]), .B1(n_0_0_72), .B2(multiplier[30]), .ZN(
      n_0_0_50));
   OAI221_X1 i_0_0_183 (.A(n_0_0_52), .B1(n_0_0_55), .B2(n_0_0_75), .C1(
      multiplier[22]), .C2(n_0_0_72), .ZN(n_0_0_51));
   AOI21_X1 i_0_0_184 (.A(n_0_0_53), .B1(n_0_0_56), .B2(n_0_0_57), .ZN(n_0_0_52));
   OAI22_X1 i_0_0_185 (.A1(n_0_0_74), .A2(n_0_0_54), .B1(n_0_0_70), .B2(
      multiplier[23]), .ZN(n_0_0_53));
   MUX2_X1 i_0_0_186 (.A(multiplier[18]), .B(multiplier[19]), .S(ctr[0]), 
      .Z(n_0_0_54));
   MUX2_X1 i_0_0_187 (.A(multiplier[20]), .B(multiplier[21]), .S(ctr[0]), 
      .Z(n_0_0_55));
   AOI21_X1 i_0_0_188 (.A(n_0_0_76), .B1(multiplier[17]), .B2(ctr[0]), .ZN(
      n_0_0_56));
   NAND2_X1 i_0_0_189 (.A1(n_0_0_117), .A2(multiplier[16]), .ZN(n_0_0_57));
   OAI33_X1 i_0_0_190 (.A1(n_0_0_65), .A2(n_0_0_69), .A3(n_0_0_66), .B1(n_0_0_60), 
      .B2(n_0_0_59), .B3(ctr[3]), .ZN(n_0_0_58));
   OAI221_X1 i_0_0_191 (.A(n_0_0_62), .B1(multiplier[7]), .B2(n_0_0_70), 
      .C1(n_0_0_64), .C2(n_0_0_76), .ZN(n_0_0_59));
   OAI22_X1 i_0_0_192 (.A1(n_0_0_74), .A2(n_0_0_61), .B1(n_0_0_72), .B2(
      multiplier[6]), .ZN(n_0_0_60));
   MUX2_X1 i_0_0_193 (.A(multiplier[2]), .B(multiplier[3]), .S(ctr[0]), .Z(
      n_0_0_61));
   OAI21_X1 i_0_0_194 (.A(n_0_0_63), .B1(n_0_0_114), .B2(ctr[0]), .ZN(n_0_0_62));
   AOI21_X1 i_0_0_195 (.A(n_0_0_75), .B1(multiplier[5]), .B2(ctr[0]), .ZN(
      n_0_0_63));
   MUX2_X1 i_0_0_196 (.A(multiplier[0]), .B(multiplier[1]), .S(ctr[0]), .Z(
      n_0_0_64));
   OAI221_X1 i_0_0_197 (.A(n_0_0_67), .B1(n_0_0_71), .B2(n_0_0_75), .C1(
      multiplier[14]), .C2(n_0_0_72), .ZN(n_0_0_65));
   OAI21_X1 i_0_0_198 (.A(ctr[3]), .B1(n_0_0_76), .B2(n_0_0_73), .ZN(n_0_0_66));
   OAI21_X1 i_0_0_199 (.A(n_0_0_68), .B1(n_0_0_115), .B2(ctr[0]), .ZN(n_0_0_67));
   AOI21_X1 i_0_0_200 (.A(n_0_0_74), .B1(multiplier[11]), .B2(ctr[0]), .ZN(
      n_0_0_68));
   NOR2_X1 i_0_0_201 (.A1(n_0_0_70), .A2(multiplier[15]), .ZN(n_0_0_69));
   NAND3_X1 i_0_0_202 (.A1(ctr[2]), .A2(ctr[1]), .A3(ctr[0]), .ZN(n_0_0_70));
   MUX2_X1 i_0_0_203 (.A(multiplier[12]), .B(multiplier[13]), .S(ctr[0]), 
      .Z(n_0_0_71));
   NAND3_X1 i_0_0_204 (.A1(n_0_0_117), .A2(ctr[1]), .A3(ctr[2]), .ZN(n_0_0_72));
   MUX2_X1 i_0_0_205 (.A(multiplier[8]), .B(multiplier[9]), .S(ctr[0]), .Z(
      n_0_0_73));
   OR2_X1 i_0_0_206 (.A1(n_0_0_118), .A2(ctr[2]), .ZN(n_0_0_74));
   NAND2_X1 i_0_0_207 (.A1(n_0_0_118), .A2(ctr[2]), .ZN(n_0_0_75));
   OR2_X1 i_0_0_208 (.A1(ctr[2]), .A2(ctr[1]), .ZN(n_0_0_76));
   MUX2_X1 i_0_0_209 (.A(n_0_13), .B(n_0_340), .S(n_0_0_77), .Z(n_0_276));
   MUX2_X1 i_0_0_210 (.A(n_0_14), .B(n_0_341), .S(n_0_0_77), .Z(n_0_277));
   MUX2_X1 i_0_0_211 (.A(n_0_15), .B(n_0_342), .S(n_0_0_77), .Z(n_0_278));
   MUX2_X1 i_0_0_212 (.A(n_0_16), .B(n_0_343), .S(n_0_0_77), .Z(n_0_279));
   MUX2_X1 i_0_0_213 (.A(n_0_17), .B(n_0_344), .S(n_0_0_77), .Z(n_0_280));
   MUX2_X1 i_0_0_214 (.A(n_0_18), .B(n_0_345), .S(n_0_0_77), .Z(n_0_281));
   MUX2_X1 i_0_0_215 (.A(n_0_19), .B(n_0_346), .S(n_0_0_77), .Z(n_0_282));
   MUX2_X1 i_0_0_216 (.A(n_0_20), .B(n_0_347), .S(n_0_0_77), .Z(n_0_283));
   MUX2_X1 i_0_0_217 (.A(n_0_21), .B(n_0_348), .S(n_0_0_77), .Z(n_0_284));
   MUX2_X1 i_0_0_218 (.A(n_0_22), .B(n_0_349), .S(n_0_0_77), .Z(n_0_285));
   MUX2_X1 i_0_0_219 (.A(n_0_23), .B(n_0_350), .S(n_0_0_77), .Z(n_0_286));
   MUX2_X1 i_0_0_220 (.A(n_0_24), .B(n_0_351), .S(n_0_0_77), .Z(n_0_287));
   MUX2_X1 i_0_0_221 (.A(n_0_25), .B(n_0_352), .S(n_0_0_77), .Z(n_0_288));
   MUX2_X1 i_0_0_222 (.A(n_0_26), .B(n_0_353), .S(n_0_0_77), .Z(n_0_289));
   MUX2_X1 i_0_0_223 (.A(n_0_27), .B(n_0_354), .S(n_0_0_77), .Z(n_0_290));
   MUX2_X1 i_0_0_224 (.A(n_0_28), .B(n_0_355), .S(n_0_0_77), .Z(n_0_291));
   MUX2_X1 i_0_0_225 (.A(n_0_29), .B(n_0_356), .S(n_0_0_77), .Z(n_0_292));
   MUX2_X1 i_0_0_226 (.A(n_0_30), .B(n_0_357), .S(n_0_0_77), .Z(n_0_293));
   MUX2_X1 i_0_0_227 (.A(n_0_31), .B(n_0_358), .S(n_0_0_77), .Z(n_0_294));
   MUX2_X1 i_0_0_228 (.A(n_0_32), .B(n_0_359), .S(n_0_0_77), .Z(n_0_295));
   MUX2_X1 i_0_0_229 (.A(n_0_33), .B(n_0_360), .S(n_0_0_77), .Z(n_0_296));
   MUX2_X1 i_0_0_230 (.A(n_0_34), .B(n_0_361), .S(n_0_0_77), .Z(n_0_297));
   MUX2_X1 i_0_0_231 (.A(n_0_35), .B(n_0_362), .S(n_0_0_77), .Z(n_0_298));
   MUX2_X1 i_0_0_232 (.A(n_0_36), .B(n_0_363), .S(n_0_0_77), .Z(n_0_299));
   MUX2_X1 i_0_0_233 (.A(n_0_37), .B(n_0_364), .S(n_0_0_77), .Z(n_0_300));
   MUX2_X1 i_0_0_234 (.A(n_0_38), .B(n_0_365), .S(n_0_0_77), .Z(n_0_301));
   MUX2_X1 i_0_0_235 (.A(n_0_39), .B(n_0_366), .S(n_0_0_77), .Z(n_0_302));
   MUX2_X1 i_0_0_236 (.A(n_0_40), .B(n_0_367), .S(n_0_0_77), .Z(n_0_303));
   MUX2_X1 i_0_0_237 (.A(n_0_41), .B(n_0_368), .S(n_0_0_77), .Z(n_0_304));
   MUX2_X1 i_0_0_238 (.A(n_0_42), .B(n_0_369), .S(n_0_0_77), .Z(n_0_305));
   NAND2_X1 i_0_0_239 (.A1(rst), .A2(n_0_370), .ZN(n_0_0_77));
   NOR2_X1 i_0_0_240 (.A1(n_0_0_119), .A2(n_0_0_79), .ZN(n_0_0_78));
   AOI21_X1 i_0_0_241 (.A(n_0_0_79), .B1(n_0_0_116), .B2(rst), .ZN(n_0_306));
   MUX2_X1 i_0_0_242 (.A(y[0]), .B(x[0]), .S(x[31]), .Z(n_0_307));
   MUX2_X1 i_0_0_243 (.A(y[1]), .B(x[1]), .S(x[31]), .Z(n_0_308));
   MUX2_X1 i_0_0_244 (.A(y[2]), .B(x[2]), .S(x[31]), .Z(n_0_309));
   MUX2_X1 i_0_0_245 (.A(y[3]), .B(x[3]), .S(x[31]), .Z(n_0_310));
   MUX2_X1 i_0_0_246 (.A(y[4]), .B(x[4]), .S(x[31]), .Z(n_0_311));
   MUX2_X1 i_0_0_247 (.A(y[5]), .B(x[5]), .S(x[31]), .Z(n_0_312));
   MUX2_X1 i_0_0_248 (.A(y[6]), .B(x[6]), .S(x[31]), .Z(n_0_313));
   MUX2_X1 i_0_0_249 (.A(y[7]), .B(x[7]), .S(x[31]), .Z(n_0_314));
   MUX2_X1 i_0_0_250 (.A(y[8]), .B(x[8]), .S(x[31]), .Z(n_0_315));
   MUX2_X1 i_0_0_251 (.A(y[9]), .B(x[9]), .S(x[31]), .Z(n_0_316));
   MUX2_X1 i_0_0_252 (.A(y[10]), .B(x[10]), .S(x[31]), .Z(n_0_317));
   MUX2_X1 i_0_0_253 (.A(y[11]), .B(x[11]), .S(x[31]), .Z(n_0_318));
   MUX2_X1 i_0_0_254 (.A(y[12]), .B(x[12]), .S(x[31]), .Z(n_0_319));
   MUX2_X1 i_0_0_255 (.A(y[13]), .B(x[13]), .S(x[31]), .Z(n_0_320));
   MUX2_X1 i_0_0_256 (.A(y[14]), .B(x[14]), .S(x[31]), .Z(n_0_321));
   MUX2_X1 i_0_0_257 (.A(y[15]), .B(x[15]), .S(x[31]), .Z(n_0_322));
   MUX2_X1 i_0_0_258 (.A(y[16]), .B(x[16]), .S(x[31]), .Z(n_0_323));
   MUX2_X1 i_0_0_259 (.A(y[17]), .B(x[17]), .S(x[31]), .Z(n_0_324));
   MUX2_X1 i_0_0_260 (.A(y[18]), .B(x[18]), .S(x[31]), .Z(n_0_325));
   MUX2_X1 i_0_0_261 (.A(y[19]), .B(x[19]), .S(x[31]), .Z(n_0_326));
   MUX2_X1 i_0_0_262 (.A(y[20]), .B(x[20]), .S(x[31]), .Z(n_0_327));
   MUX2_X1 i_0_0_263 (.A(y[21]), .B(x[21]), .S(x[31]), .Z(n_0_328));
   MUX2_X1 i_0_0_264 (.A(y[22]), .B(x[22]), .S(x[31]), .Z(n_0_329));
   MUX2_X1 i_0_0_265 (.A(y[23]), .B(x[23]), .S(x[31]), .Z(n_0_330));
   MUX2_X1 i_0_0_266 (.A(y[24]), .B(x[24]), .S(x[31]), .Z(n_0_331));
   MUX2_X1 i_0_0_267 (.A(y[25]), .B(x[25]), .S(x[31]), .Z(n_0_332));
   MUX2_X1 i_0_0_268 (.A(y[26]), .B(x[26]), .S(x[31]), .Z(n_0_333));
   MUX2_X1 i_0_0_269 (.A(y[27]), .B(x[27]), .S(x[31]), .Z(n_0_334));
   MUX2_X1 i_0_0_270 (.A(y[28]), .B(x[28]), .S(x[31]), .Z(n_0_335));
   MUX2_X1 i_0_0_271 (.A(y[29]), .B(x[29]), .S(x[31]), .Z(n_0_336));
   MUX2_X1 i_0_0_272 (.A(y[30]), .B(x[30]), .S(x[31]), .Z(n_0_337));
   OR2_X1 i_0_0_273 (.A1(x[31]), .A2(y[31]), .ZN(n_0_338));
   MUX2_X1 i_0_0_274 (.A(x[0]), .B(y[0]), .S(x[31]), .Z(n_0_339));
   MUX2_X1 i_0_0_275 (.A(x[1]), .B(y[1]), .S(x[31]), .Z(n_0_340));
   MUX2_X1 i_0_0_276 (.A(x[2]), .B(y[2]), .S(x[31]), .Z(n_0_341));
   MUX2_X1 i_0_0_277 (.A(x[3]), .B(y[3]), .S(x[31]), .Z(n_0_342));
   MUX2_X1 i_0_0_278 (.A(x[4]), .B(y[4]), .S(x[31]), .Z(n_0_343));
   MUX2_X1 i_0_0_279 (.A(x[5]), .B(y[5]), .S(x[31]), .Z(n_0_344));
   MUX2_X1 i_0_0_280 (.A(x[6]), .B(y[6]), .S(x[31]), .Z(n_0_345));
   MUX2_X1 i_0_0_281 (.A(x[7]), .B(y[7]), .S(x[31]), .Z(n_0_346));
   MUX2_X1 i_0_0_282 (.A(x[8]), .B(y[8]), .S(x[31]), .Z(n_0_347));
   MUX2_X1 i_0_0_283 (.A(x[9]), .B(y[9]), .S(x[31]), .Z(n_0_348));
   MUX2_X1 i_0_0_284 (.A(x[10]), .B(y[10]), .S(x[31]), .Z(n_0_349));
   MUX2_X1 i_0_0_285 (.A(x[11]), .B(y[11]), .S(x[31]), .Z(n_0_350));
   MUX2_X1 i_0_0_286 (.A(x[12]), .B(y[12]), .S(x[31]), .Z(n_0_351));
   MUX2_X1 i_0_0_287 (.A(x[13]), .B(y[13]), .S(x[31]), .Z(n_0_352));
   MUX2_X1 i_0_0_288 (.A(x[14]), .B(y[14]), .S(x[31]), .Z(n_0_353));
   MUX2_X1 i_0_0_289 (.A(x[15]), .B(y[15]), .S(x[31]), .Z(n_0_354));
   MUX2_X1 i_0_0_290 (.A(x[16]), .B(y[16]), .S(x[31]), .Z(n_0_355));
   MUX2_X1 i_0_0_291 (.A(x[17]), .B(y[17]), .S(x[31]), .Z(n_0_356));
   MUX2_X1 i_0_0_292 (.A(x[18]), .B(y[18]), .S(x[31]), .Z(n_0_357));
   MUX2_X1 i_0_0_293 (.A(x[19]), .B(y[19]), .S(x[31]), .Z(n_0_358));
   MUX2_X1 i_0_0_294 (.A(x[20]), .B(y[20]), .S(x[31]), .Z(n_0_359));
   MUX2_X1 i_0_0_295 (.A(x[21]), .B(y[21]), .S(x[31]), .Z(n_0_360));
   MUX2_X1 i_0_0_296 (.A(x[22]), .B(y[22]), .S(x[31]), .Z(n_0_361));
   MUX2_X1 i_0_0_297 (.A(x[23]), .B(y[23]), .S(x[31]), .Z(n_0_362));
   MUX2_X1 i_0_0_298 (.A(x[24]), .B(y[24]), .S(x[31]), .Z(n_0_363));
   MUX2_X1 i_0_0_299 (.A(x[25]), .B(y[25]), .S(x[31]), .Z(n_0_364));
   MUX2_X1 i_0_0_300 (.A(x[26]), .B(y[26]), .S(x[31]), .Z(n_0_365));
   MUX2_X1 i_0_0_301 (.A(x[27]), .B(y[27]), .S(x[31]), .Z(n_0_366));
   MUX2_X1 i_0_0_302 (.A(x[28]), .B(y[28]), .S(x[31]), .Z(n_0_367));
   MUX2_X1 i_0_0_303 (.A(x[29]), .B(y[29]), .S(x[31]), .Z(n_0_368));
   MUX2_X1 i_0_0_304 (.A(x[30]), .B(y[30]), .S(x[31]), .Z(n_0_369));
   INV_X1 i_0_0_305 (.A(n_0_0_79), .ZN(n_0_370));
   NAND2_X1 i_0_0_306 (.A1(x[31]), .A2(y[31]), .ZN(n_0_0_79));
   INV_X1 i_0_0_307 (.A(n_0_0_80), .ZN(n_0_371));
   NOR2_X1 i_0_0_308 (.A1(rst), .A2(ctr[5]), .ZN(n_0_0_80));
   INV_X1 i_0_0_309 (.A(n_0_74), .ZN(n_0_0_81));
   INV_X1 i_0_0_310 (.A(n_0_459), .ZN(n_0_0_82));
   INV_X1 i_0_0_311 (.A(n_0_458), .ZN(n_0_0_83));
   INV_X1 i_0_0_312 (.A(n_0_457), .ZN(n_0_0_84));
   INV_X1 i_0_0_313 (.A(n_0_456), .ZN(n_0_0_85));
   INV_X1 i_0_0_314 (.A(n_0_455), .ZN(n_0_0_86));
   INV_X1 i_0_0_315 (.A(n_0_454), .ZN(n_0_0_87));
   INV_X1 i_0_0_316 (.A(n_0_453), .ZN(n_0_0_88));
   INV_X1 i_0_0_317 (.A(n_0_452), .ZN(n_0_0_89));
   INV_X1 i_0_0_318 (.A(n_0_451), .ZN(n_0_0_90));
   INV_X1 i_0_0_319 (.A(n_0_450), .ZN(n_0_0_91));
   INV_X1 i_0_0_320 (.A(n_0_449), .ZN(n_0_0_92));
   INV_X1 i_0_0_321 (.A(n_0_448), .ZN(n_0_0_93));
   INV_X1 i_0_0_322 (.A(n_0_447), .ZN(n_0_0_94));
   INV_X1 i_0_0_323 (.A(n_0_446), .ZN(n_0_0_95));
   INV_X1 i_0_0_324 (.A(n_0_445), .ZN(n_0_0_96));
   INV_X1 i_0_0_325 (.A(n_0_444), .ZN(n_0_0_97));
   INV_X1 i_0_0_326 (.A(n_0_443), .ZN(n_0_0_98));
   INV_X1 i_0_0_327 (.A(n_0_442), .ZN(n_0_0_99));
   INV_X1 i_0_0_328 (.A(n_0_441), .ZN(n_0_0_100));
   INV_X1 i_0_0_329 (.A(n_0_440), .ZN(n_0_0_101));
   INV_X1 i_0_0_330 (.A(n_0_439), .ZN(n_0_0_102));
   INV_X1 i_0_0_331 (.A(n_0_438), .ZN(n_0_0_103));
   INV_X1 i_0_0_332 (.A(n_0_437), .ZN(n_0_0_104));
   INV_X1 i_0_0_333 (.A(n_0_436), .ZN(n_0_0_105));
   INV_X1 i_0_0_334 (.A(n_0_435), .ZN(n_0_0_106));
   INV_X1 i_0_0_335 (.A(n_0_434), .ZN(n_0_0_107));
   INV_X1 i_0_0_336 (.A(n_0_433), .ZN(n_0_0_108));
   INV_X1 i_0_0_337 (.A(n_0_432), .ZN(n_0_0_109));
   INV_X1 i_0_0_338 (.A(n_0_431), .ZN(n_0_0_110));
   INV_X1 i_0_0_339 (.A(n_0_430), .ZN(n_0_0_111));
   INV_X1 i_0_0_340 (.A(n_0_429), .ZN(n_0_0_112));
   INV_X1 i_0_0_341 (.A(n_0_428), .ZN(n_0_0_113));
   INV_X1 i_0_0_342 (.A(multiplier[4]), .ZN(n_0_0_114));
   INV_X1 i_0_0_343 (.A(multiplier[10]), .ZN(n_0_0_115));
   INV_X1 i_0_0_344 (.A(n_0_43), .ZN(n_0_0_116));
   INV_X1 i_0_0_345 (.A(ctr[0]), .ZN(n_0_0_117));
   INV_X1 i_0_0_346 (.A(ctr[1]), .ZN(n_0_0_118));
   INV_X1 i_0_0_347 (.A(rst), .ZN(n_0_0_119));
   DFF_X1 \multiplicand_reg[63]  (.D(n_0_273), .CK(n_0_373), .Q(n_0_372), .QN());
   DFF_X1 \multiplicand_reg[62]  (.D(n_0_272), .CK(n_0_373), .Q(n_0_428), .QN());
   DFF_X1 \multiplicand_reg[61]  (.D(n_0_271), .CK(n_0_373), .Q(n_0_429), .QN());
   DFF_X1 \multiplicand_reg[60]  (.D(n_0_270), .CK(n_0_373), .Q(n_0_430), .QN());
   DFF_X1 \multiplicand_reg[59]  (.D(n_0_269), .CK(n_0_373), .Q(n_0_431), .QN());
   DFF_X1 \multiplicand_reg[58]  (.D(n_0_268), .CK(n_0_373), .Q(n_0_432), .QN());
   DFF_X1 \multiplicand_reg[57]  (.D(n_0_267), .CK(n_0_373), .Q(n_0_433), .QN());
   DFF_X1 \multiplicand_reg[56]  (.D(n_0_266), .CK(n_0_373), .Q(n_0_434), .QN());
   DFF_X1 \multiplicand_reg[55]  (.D(n_0_265), .CK(n_0_373), .Q(n_0_435), .QN());
   DFF_X1 \multiplicand_reg[54]  (.D(n_0_264), .CK(n_0_373), .Q(n_0_436), .QN());
   DFF_X1 \multiplicand_reg[53]  (.D(n_0_263), .CK(n_0_373), .Q(n_0_437), .QN());
   DFF_X1 \multiplicand_reg[52]  (.D(n_0_262), .CK(n_0_373), .Q(n_0_438), .QN());
   DFF_X1 \multiplicand_reg[51]  (.D(n_0_261), .CK(n_0_373), .Q(n_0_439), .QN());
   DFF_X1 \multiplicand_reg[50]  (.D(n_0_260), .CK(n_0_373), .Q(n_0_440), .QN());
   DFF_X1 \multiplicand_reg[49]  (.D(n_0_259), .CK(n_0_373), .Q(n_0_441), .QN());
   DFF_X1 \multiplicand_reg[48]  (.D(n_0_258), .CK(n_0_373), .Q(n_0_442), .QN());
   DFF_X1 \multiplicand_reg[47]  (.D(n_0_257), .CK(n_0_373), .Q(n_0_443), .QN());
   DFF_X1 \multiplicand_reg[46]  (.D(n_0_256), .CK(n_0_373), .Q(n_0_444), .QN());
   DFF_X1 \multiplicand_reg[45]  (.D(n_0_255), .CK(n_0_373), .Q(n_0_445), .QN());
   DFF_X1 \multiplicand_reg[44]  (.D(n_0_254), .CK(n_0_373), .Q(n_0_446), .QN());
   DFF_X1 \multiplicand_reg[43]  (.D(n_0_253), .CK(n_0_373), .Q(n_0_447), .QN());
   DFF_X1 \multiplicand_reg[42]  (.D(n_0_252), .CK(n_0_373), .Q(n_0_448), .QN());
   DFF_X1 \multiplicand_reg[41]  (.D(n_0_251), .CK(n_0_373), .Q(n_0_449), .QN());
   DFF_X1 \multiplicand_reg[40]  (.D(n_0_250), .CK(n_0_373), .Q(n_0_450), .QN());
   DFF_X1 \multiplicand_reg[39]  (.D(n_0_249), .CK(n_0_373), .Q(n_0_451), .QN());
   DFF_X1 \multiplicand_reg[38]  (.D(n_0_248), .CK(n_0_373), .Q(n_0_452), .QN());
   DFF_X1 \multiplicand_reg[37]  (.D(n_0_247), .CK(n_0_373), .Q(n_0_453), .QN());
   DFF_X1 \multiplicand_reg[36]  (.D(n_0_246), .CK(n_0_373), .Q(n_0_454), .QN());
   DFF_X1 \multiplicand_reg[35]  (.D(n_0_245), .CK(n_0_373), .Q(n_0_455), .QN());
   DFF_X1 \multiplicand_reg[34]  (.D(n_0_244), .CK(n_0_373), .Q(n_0_456), .QN());
   DFF_X1 \multiplicand_reg[33]  (.D(n_0_243), .CK(n_0_373), .Q(n_0_457), .QN());
   DFF_X1 \multiplicand_reg[32]  (.D(n_0_242), .CK(n_0_373), .Q(n_0_458), .QN());
   DFF_X1 \multiplicand_reg[31]  (.D(n_0_241), .CK(n_0_373), .Q(n_0_459), .QN());
   DFF_X1 \multiplicand_reg[30]  (.D(n_0_240), .CK(n_0_373), .Q(n_0_460), .QN());
   DFF_X1 \multiplicand_reg[29]  (.D(n_0_239), .CK(n_0_373), .Q(n_0_461), .QN());
   DFF_X1 \multiplicand_reg[28]  (.D(n_0_238), .CK(n_0_373), .Q(n_0_462), .QN());
   DFF_X1 \multiplicand_reg[27]  (.D(n_0_237), .CK(n_0_373), .Q(n_0_463), .QN());
   DFF_X1 \multiplicand_reg[26]  (.D(n_0_236), .CK(n_0_373), .Q(n_0_464), .QN());
   DFF_X1 \multiplicand_reg[25]  (.D(n_0_235), .CK(n_0_373), .Q(n_0_465), .QN());
   DFF_X1 \multiplicand_reg[24]  (.D(n_0_234), .CK(n_0_373), .Q(n_0_466), .QN());
   DFF_X1 \multiplicand_reg[23]  (.D(n_0_233), .CK(n_0_373), .Q(n_0_467), .QN());
   DFF_X1 \multiplicand_reg[22]  (.D(n_0_232), .CK(n_0_373), .Q(n_0_468), .QN());
   DFF_X1 \multiplicand_reg[21]  (.D(n_0_231), .CK(n_0_373), .Q(n_0_469), .QN());
   DFF_X1 \multiplicand_reg[20]  (.D(n_0_230), .CK(n_0_373), .Q(n_0_470), .QN());
   DFF_X1 \multiplicand_reg[19]  (.D(n_0_229), .CK(n_0_373), .Q(n_0_471), .QN());
   DFF_X1 \multiplicand_reg[18]  (.D(n_0_228), .CK(n_0_373), .Q(n_0_472), .QN());
   DFF_X1 \multiplicand_reg[17]  (.D(n_0_227), .CK(n_0_373), .Q(n_0_473), .QN());
   DFF_X1 \multiplicand_reg[16]  (.D(n_0_226), .CK(n_0_373), .Q(n_0_474), .QN());
   DFF_X1 \multiplicand_reg[15]  (.D(n_0_225), .CK(n_0_373), .Q(n_0_475), .QN());
   DFF_X1 \multiplicand_reg[14]  (.D(n_0_224), .CK(n_0_373), .Q(n_0_476), .QN());
   DFF_X1 \multiplicand_reg[13]  (.D(n_0_223), .CK(n_0_373), .Q(n_0_477), .QN());
   DFF_X1 \multiplicand_reg[12]  (.D(n_0_222), .CK(n_0_373), .Q(n_0_478), .QN());
   DFF_X1 \multiplicand_reg[11]  (.D(n_0_221), .CK(n_0_373), .Q(n_0_479), .QN());
   DFF_X1 \multiplicand_reg[10]  (.D(n_0_220), .CK(n_0_373), .Q(n_0_480), .QN());
   DFF_X1 \multiplicand_reg[9]  (.D(n_0_219), .CK(n_0_373), .Q(n_0_481), .QN());
   DFF_X1 \multiplicand_reg[8]  (.D(n_0_218), .CK(n_0_373), .Q(n_0_482), .QN());
   DFF_X1 \multiplicand_reg[7]  (.D(n_0_217), .CK(n_0_373), .Q(n_0_483), .QN());
   DFF_X1 \multiplicand_reg[6]  (.D(n_0_216), .CK(n_0_373), .Q(n_0_484), .QN());
   DFF_X1 \multiplicand_reg[5]  (.D(n_0_215), .CK(n_0_373), .Q(n_0_485), .QN());
   DFF_X1 \multiplicand_reg[4]  (.D(n_0_214), .CK(n_0_373), .Q(n_0_486), .QN());
   DFF_X1 \multiplicand_reg[3]  (.D(n_0_213), .CK(n_0_373), .Q(n_0_487), .QN());
   DFF_X1 \multiplicand_reg[2]  (.D(n_0_212), .CK(n_0_373), .Q(n_0_488), .QN());
   DFF_X1 \multiplicand_reg[1]  (.D(n_0_211), .CK(n_0_373), .Q(n_0_489), .QN());
   DFF_X1 \multiplicand_reg[0]  (.D(n_0_210), .CK(n_0_373), .Q(n_0_490), .QN());
   CLKGATETST_X1 clk_gate_accumulator_reg (.CK(clk), .E(n_0_275), .SE(1'b0), 
      .GCK(n_0_374));
   DFF_X1 \accumulator_reg[63]  (.D(n_0_203), .CK(n_0_374), .Q(n_0_375), .QN());
   DFF_X1 \accumulator_reg[62]  (.D(n_0_202), .CK(n_0_374), .Q(n_0_376), .QN());
   DFF_X1 \accumulator_reg[61]  (.D(n_0_201), .CK(n_0_374), .Q(n_0_377), .QN());
   DFF_X1 \accumulator_reg[60]  (.D(n_0_200), .CK(n_0_374), .Q(n_0_378), .QN());
   DFF_X1 \accumulator_reg[59]  (.D(n_0_199), .CK(n_0_374), .Q(n_0_379), .QN());
   DFF_X1 \accumulator_reg[58]  (.D(n_0_198), .CK(n_0_374), .Q(n_0_380), .QN());
   DFF_X1 \accumulator_reg[57]  (.D(n_0_197), .CK(n_0_374), .Q(n_0_381), .QN());
   DFF_X1 \accumulator_reg[56]  (.D(n_0_196), .CK(n_0_374), .Q(n_0_382), .QN());
   DFF_X1 \accumulator_reg[55]  (.D(n_0_195), .CK(n_0_374), .Q(n_0_383), .QN());
   DFF_X1 \accumulator_reg[54]  (.D(n_0_194), .CK(n_0_374), .Q(n_0_384), .QN());
   DFF_X1 \accumulator_reg[53]  (.D(n_0_193), .CK(n_0_374), .Q(n_0_385), .QN());
   DFF_X1 \accumulator_reg[52]  (.D(n_0_192), .CK(n_0_374), .Q(n_0_386), .QN());
   DFF_X1 \accumulator_reg[51]  (.D(n_0_191), .CK(n_0_374), .Q(n_0_387), .QN());
   DFF_X1 \accumulator_reg[50]  (.D(n_0_190), .CK(n_0_374), .Q(n_0_388), .QN());
   DFF_X1 \accumulator_reg[49]  (.D(n_0_189), .CK(n_0_374), .Q(n_0_389), .QN());
   DFF_X1 \accumulator_reg[48]  (.D(n_0_188), .CK(n_0_374), .Q(n_0_390), .QN());
   DFF_X1 \accumulator_reg[47]  (.D(n_0_187), .CK(n_0_374), .Q(n_0_391), .QN());
   DFF_X1 \accumulator_reg[46]  (.D(n_0_186), .CK(n_0_374), .Q(n_0_392), .QN());
   DFF_X1 \accumulator_reg[45]  (.D(n_0_185), .CK(n_0_374), .Q(n_0_393), .QN());
   DFF_X1 \accumulator_reg[44]  (.D(n_0_184), .CK(n_0_374), .Q(n_0_394), .QN());
   DFF_X1 \accumulator_reg[43]  (.D(n_0_183), .CK(n_0_374), .Q(n_0_395), .QN());
   DFF_X1 \accumulator_reg[42]  (.D(n_0_182), .CK(n_0_374), .Q(n_0_396), .QN());
   DFF_X1 \accumulator_reg[41]  (.D(n_0_181), .CK(n_0_374), .Q(n_0_397), .QN());
   DFF_X1 \accumulator_reg[40]  (.D(n_0_180), .CK(n_0_374), .Q(n_0_398), .QN());
   DFF_X1 \accumulator_reg[39]  (.D(n_0_179), .CK(n_0_374), .Q(n_0_399), .QN());
   DFF_X1 \accumulator_reg[38]  (.D(n_0_178), .CK(n_0_374), .Q(n_0_400), .QN());
   DFF_X1 \accumulator_reg[37]  (.D(n_0_177), .CK(n_0_374), .Q(n_0_401), .QN());
   DFF_X1 \accumulator_reg[36]  (.D(n_0_176), .CK(n_0_374), .Q(n_0_402), .QN());
   DFF_X1 \accumulator_reg[35]  (.D(n_0_175), .CK(n_0_374), .Q(n_0_403), .QN());
   DFF_X1 \accumulator_reg[34]  (.D(n_0_174), .CK(n_0_374), .Q(n_0_404), .QN());
   DFF_X1 \accumulator_reg[33]  (.D(n_0_173), .CK(n_0_374), .Q(n_0_405), .QN());
   DFF_X1 \accumulator_reg[32]  (.D(n_0_172), .CK(n_0_374), .Q(n_0_406), .QN());
   DFF_X1 \accumulator_reg[31]  (.D(n_0_171), .CK(n_0_374), .Q(n_0_407), .QN());
   DFF_X1 \accumulator_reg[30]  (.D(n_0_170), .CK(n_0_374), .Q(n_0_408), .QN());
   DFF_X1 \accumulator_reg[29]  (.D(n_0_169), .CK(n_0_374), .Q(n_0_409), .QN());
   DFF_X1 \accumulator_reg[28]  (.D(n_0_168), .CK(n_0_374), .Q(n_0_410), .QN());
   DFF_X1 \accumulator_reg[27]  (.D(n_0_167), .CK(n_0_374), .Q(n_0_411), .QN());
   DFF_X1 \accumulator_reg[26]  (.D(n_0_166), .CK(n_0_374), .Q(n_0_412), .QN());
   DFF_X1 \accumulator_reg[25]  (.D(n_0_165), .CK(n_0_374), .Q(n_0_413), .QN());
   DFF_X1 \accumulator_reg[24]  (.D(n_0_164), .CK(n_0_374), .Q(n_0_414), .QN());
   DFF_X1 \accumulator_reg[23]  (.D(n_0_163), .CK(n_0_374), .Q(n_0_415), .QN());
   DFF_X1 \accumulator_reg[22]  (.D(n_0_162), .CK(n_0_374), .Q(n_0_416), .QN());
   DFF_X1 \accumulator_reg[21]  (.D(n_0_161), .CK(n_0_374), .Q(n_0_417), .QN());
   DFF_X1 \accumulator_reg[20]  (.D(n_0_160), .CK(n_0_374), .Q(n_0_418), .QN());
   DFF_X1 \accumulator_reg[19]  (.D(n_0_159), .CK(n_0_374), .Q(n_0_419), .QN());
   DFF_X1 \accumulator_reg[18]  (.D(n_0_158), .CK(n_0_374), .Q(n_0_420), .QN());
   DFF_X1 \accumulator_reg[17]  (.D(n_0_157), .CK(n_0_374), .Q(n_0_421), .QN());
   DFF_X1 \accumulator_reg[16]  (.D(n_0_156), .CK(n_0_374), .Q(n_0_422), .QN());
   DFF_X1 \accumulator_reg[15]  (.D(n_0_155), .CK(n_0_374), .Q(n_0_423), .QN());
   DFF_X1 \accumulator_reg[14]  (.D(n_0_154), .CK(n_0_374), .Q(n_0_424), .QN());
   DFF_X1 \accumulator_reg[13]  (.D(n_0_153), .CK(n_0_374), .Q(n_0_425), .QN());
   DFF_X1 \accumulator_reg[12]  (.D(n_0_152), .CK(n_0_374), .Q(n_0_426), .QN());
   DFF_X1 \accumulator_reg[11]  (.D(n_0_151), .CK(n_0_374), .Q(n_0_427), .QN());
   DFF_X1 \accumulator_reg[10]  (.D(n_0_150), .CK(n_0_374), .Q(n_0_1), .QN());
   DFF_X1 \accumulator_reg[9]  (.D(n_0_149), .CK(n_0_374), .Q(n_0_2), .QN());
   DFF_X1 \accumulator_reg[8]  (.D(n_0_148), .CK(n_0_374), .Q(n_0_3), .QN());
   DFF_X1 \accumulator_reg[7]  (.D(n_0_147), .CK(n_0_374), .Q(n_0_4), .QN());
   DFF_X1 \accumulator_reg[6]  (.D(n_0_146), .CK(n_0_374), .Q(n_0_5), .QN());
   DFF_X1 \accumulator_reg[5]  (.D(n_0_145), .CK(n_0_374), .Q(n_0_6), .QN());
   DFF_X1 \accumulator_reg[4]  (.D(n_0_144), .CK(n_0_374), .Q(n_0_7), .QN());
   DFF_X1 \accumulator_reg[3]  (.D(n_0_143), .CK(n_0_374), .Q(n_0_8), .QN());
   DFF_X1 \accumulator_reg[2]  (.D(n_0_142), .CK(n_0_374), .Q(n_0_9), .QN());
   DFF_X1 \accumulator_reg[1]  (.D(n_0_141), .CK(n_0_374), .Q(n_0_10), .QN());
   DFF_X1 \accumulator_reg[0]  (.D(n_0_140), .CK(n_0_374), .Q(n_0_11), .QN());
   CLKGATETST_X1 clk_gate_multiplier_reg (.CK(clk), .E(rst), .SE(1'b0), .GCK(
      n_0_12));
   DFF_X1 \multiplier_reg[31]  (.D(n_0_306), .CK(n_0_12), .Q(multiplier[31]), 
      .QN());
   DFF_X1 \multiplier_reg[30]  (.D(n_0_305), .CK(n_0_12), .Q(multiplier[30]), 
      .QN());
   DFF_X1 \multiplier_reg[29]  (.D(n_0_304), .CK(n_0_12), .Q(multiplier[29]), 
      .QN());
   DFF_X1 \multiplier_reg[28]  (.D(n_0_303), .CK(n_0_12), .Q(multiplier[28]), 
      .QN());
   DFF_X1 \multiplier_reg[27]  (.D(n_0_302), .CK(n_0_12), .Q(multiplier[27]), 
      .QN());
   DFF_X1 \multiplier_reg[26]  (.D(n_0_301), .CK(n_0_12), .Q(multiplier[26]), 
      .QN());
   DFF_X1 \multiplier_reg[25]  (.D(n_0_300), .CK(n_0_12), .Q(multiplier[25]), 
      .QN());
   DFF_X1 \multiplier_reg[24]  (.D(n_0_299), .CK(n_0_12), .Q(multiplier[24]), 
      .QN());
   DFF_X1 \multiplier_reg[23]  (.D(n_0_298), .CK(n_0_12), .Q(multiplier[23]), 
      .QN());
   DFF_X1 \multiplier_reg[22]  (.D(n_0_297), .CK(n_0_12), .Q(multiplier[22]), 
      .QN());
   DFF_X1 \multiplier_reg[21]  (.D(n_0_296), .CK(n_0_12), .Q(multiplier[21]), 
      .QN());
   DFF_X1 \multiplier_reg[20]  (.D(n_0_295), .CK(n_0_12), .Q(multiplier[20]), 
      .QN());
   DFF_X1 \multiplier_reg[19]  (.D(n_0_294), .CK(n_0_12), .Q(multiplier[19]), 
      .QN());
   DFF_X1 \multiplier_reg[18]  (.D(n_0_293), .CK(n_0_12), .Q(multiplier[18]), 
      .QN());
   DFF_X1 \multiplier_reg[17]  (.D(n_0_292), .CK(n_0_12), .Q(multiplier[17]), 
      .QN());
   DFF_X1 \multiplier_reg[16]  (.D(n_0_291), .CK(n_0_12), .Q(multiplier[16]), 
      .QN());
   DFF_X1 \multiplier_reg[15]  (.D(n_0_290), .CK(n_0_12), .Q(multiplier[15]), 
      .QN());
   DFF_X1 \multiplier_reg[14]  (.D(n_0_289), .CK(n_0_12), .Q(multiplier[14]), 
      .QN());
   DFF_X1 \multiplier_reg[13]  (.D(n_0_288), .CK(n_0_12), .Q(multiplier[13]), 
      .QN());
   DFF_X1 \multiplier_reg[12]  (.D(n_0_287), .CK(n_0_12), .Q(multiplier[12]), 
      .QN());
   DFF_X1 \multiplier_reg[11]  (.D(n_0_286), .CK(n_0_12), .Q(multiplier[11]), 
      .QN());
   DFF_X1 \multiplier_reg[10]  (.D(n_0_285), .CK(n_0_12), .Q(multiplier[10]), 
      .QN());
   DFF_X1 \multiplier_reg[9]  (.D(n_0_284), .CK(n_0_12), .Q(multiplier[9]), 
      .QN());
   DFF_X1 \multiplier_reg[8]  (.D(n_0_283), .CK(n_0_12), .Q(multiplier[8]), 
      .QN());
   DFF_X1 \multiplier_reg[7]  (.D(n_0_282), .CK(n_0_12), .Q(multiplier[7]), 
      .QN());
   DFF_X1 \multiplier_reg[6]  (.D(n_0_281), .CK(n_0_12), .Q(multiplier[6]), 
      .QN());
   DFF_X1 \multiplier_reg[5]  (.D(n_0_280), .CK(n_0_12), .Q(multiplier[5]), 
      .QN());
   DFF_X1 \multiplier_reg[4]  (.D(n_0_279), .CK(n_0_12), .Q(multiplier[4]), 
      .QN());
   DFF_X1 \multiplier_reg[3]  (.D(n_0_278), .CK(n_0_12), .Q(multiplier[3]), 
      .QN());
   DFF_X1 \multiplier_reg[2]  (.D(n_0_277), .CK(n_0_12), .Q(multiplier[2]), 
      .QN());
   DFF_X1 \multiplier_reg[1]  (.D(n_0_276), .CK(n_0_12), .Q(multiplier[1]), 
      .QN());
   DFF_X1 \multiplier_reg[0]  (.D(n_0_339), .CK(n_0_12), .Q(multiplier[0]), 
      .QN());
   DFF_X1 \ctr_reg[5]  (.D(n_0_209), .CK(n_0_373), .Q(ctr[5]), .QN());
   DFF_X1 \ctr_reg[4]  (.D(n_0_208), .CK(n_0_373), .Q(ctr[4]), .QN());
   DFF_X1 \ctr_reg[3]  (.D(n_0_207), .CK(n_0_373), .Q(ctr[3]), .QN());
   DFF_X1 \ctr_reg[2]  (.D(n_0_206), .CK(n_0_373), .Q(ctr[2]), .QN());
   DFF_X1 \ctr_reg[1]  (.D(n_0_205), .CK(n_0_373), .Q(ctr[1]), .QN());
   DFF_X1 \ctr_reg[0]  (.D(n_0_204), .CK(n_0_373), .Q(ctr[0]), .QN());
   CLKGATETST_X1 clk_gate_multiplicand_reg (.CK(clk), .E(n_0_274), .SE(1'b0), 
      .GCK(n_0_373));
endmodule
