
// 	Sun Jan  1 16:02:07 2023
//	vlsi
//	192.168.44.138

module registerNbits (clk_CTSPP_2, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTSPP_2;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (n_0), .D (n_33));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTSPP_2), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits

module registerNbits__2_8 (clk_CTSPP_0, clk_CTSPP_2, clk, reset, en, inp, out);

output [31:0] out;
output clk_CTSPP_0;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTSPP_2;
wire n_0_0;
wire n_1;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n6;
wire CTS_n7;
wire CTS_n8;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n8), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n8), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n8), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n7), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n7), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n7), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n7), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n7), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n7), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n7), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n7), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n7), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n7), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n7), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n7), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n7), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n8), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n8), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n8), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n8), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n8), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n8), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n8), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n8), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n8), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n8), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n8), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n8), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n8), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n8), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n8), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n8), .D (n_33));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n6), .CK (clk_CTSPP_0), .E (n_1), .SE (1'b0 ));
CLKBUF_X2 CTS_L1_c15 (.Z (clk_CTSPP_0), .A (clk_CTSPP_2));
CLKBUF_X3 CTS_L3_c5 (.Z (CTS_n7), .A (CTS_n6));
CLKBUF_X3 CTS_L3_c6 (.Z (CTS_n8), .A (CTS_n6));

endmodule //registerNbits__2_8

module registerNbits__2_5 (clk_CTSPP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTSPP_0;
wire drc_ipo_n192;
wire drc_ipo_n190;
wire drc_ipo_n188;
wire drc_ipo_n186;
wire drc_ipo_n184;
wire drc_ipo_n182;
wire drc_ipo_n180;
wire drc_ipo_n178;
wire drc_ipo_n176;
wire drc_ipo_n174;
wire drc_ipo_n172;
wire drc_ipo_n170;
wire drc_ipo_n168;
wire drc_ipo_n166;
wire drc_ipo_n164;
wire drc_ipo_n162;
wire drc_ipo_n160;
wire drc_ipo_n158;
wire drc_ipo_n156;
wire drc_ipo_n154;
wire drc_ipo_n152;
wire drc_ipo_n150;
wire drc_ipo_n148;
wire drc_ipo_n146;
wire drc_ipo_n144;
wire drc_ipo_n142;
wire drc_ipo_n140;
wire drc_ipo_n138;
wire drc_ipo_n136;
wire drc_ipo_n134;
wire drc_ipo_n132;
wire drc_ipo_n130;
wire n_0_0;
wire n_1;
wire CTS_n194;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n195;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (drc_ipo_n130), .CK (CTS_n194), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (drc_ipo_n132), .CK (CTS_n194), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (drc_ipo_n134), .CK (CTS_n194), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (drc_ipo_n136), .CK (CTS_n194), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (drc_ipo_n138), .CK (CTS_n194), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (drc_ipo_n140), .CK (CTS_n194), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (drc_ipo_n142), .CK (CTS_n194), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (drc_ipo_n144), .CK (CTS_n194), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (drc_ipo_n146), .CK (CTS_n194), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (drc_ipo_n148), .CK (CTS_n194), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (drc_ipo_n150), .CK (CTS_n194), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (drc_ipo_n152), .CK (CTS_n194), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (drc_ipo_n154), .CK (CTS_n194), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (drc_ipo_n156), .CK (CTS_n194), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (drc_ipo_n158), .CK (CTS_n194), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (drc_ipo_n160), .CK (CTS_n194), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (drc_ipo_n162), .CK (CTS_n194), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (drc_ipo_n164), .CK (CTS_n194), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (drc_ipo_n166), .CK (CTS_n194), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (drc_ipo_n168), .CK (CTS_n194), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (drc_ipo_n170), .CK (CTS_n194), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (drc_ipo_n172), .CK (CTS_n194), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (drc_ipo_n174), .CK (CTS_n194), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (drc_ipo_n176), .CK (CTS_n194), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (drc_ipo_n178), .CK (CTS_n194), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (drc_ipo_n180), .CK (CTS_n194), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (drc_ipo_n182), .CK (CTS_n194), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (drc_ipo_n184), .CK (CTS_n194), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (drc_ipo_n186), .CK (CTS_n194), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (drc_ipo_n188), .CK (CTS_n194), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (drc_ipo_n190), .CK (CTS_n194), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n192), .CK (CTS_n194), .D (n_33));
CLKGATETST_X8 clk_gate_out_reg (.GCK (CTS_n195), .CK (clk_CTSPP_0), .E (n_1), .SE (1'b0 ));
BUF_X4 drc_ipo_c96 (.Z (out[31]), .A (drc_ipo_n192));
BUF_X4 drc_ipo_c95 (.Z (out[30]), .A (drc_ipo_n190));
BUF_X4 drc_ipo_c94 (.Z (out[29]), .A (drc_ipo_n188));
CLKBUF_X2 drc_ipo_c93 (.Z (out[28]), .A (drc_ipo_n186));
BUF_X4 drc_ipo_c92 (.Z (out[27]), .A (drc_ipo_n184));
BUF_X4 drc_ipo_c91 (.Z (out[26]), .A (drc_ipo_n182));
BUF_X4 drc_ipo_c90 (.Z (out[25]), .A (drc_ipo_n180));
BUF_X4 drc_ipo_c89 (.Z (out[24]), .A (drc_ipo_n178));
BUF_X4 drc_ipo_c88 (.Z (out[23]), .A (drc_ipo_n176));
BUF_X4 drc_ipo_c87 (.Z (out[22]), .A (drc_ipo_n174));
BUF_X4 drc_ipo_c86 (.Z (out[21]), .A (drc_ipo_n172));
BUF_X4 drc_ipo_c85 (.Z (out[20]), .A (drc_ipo_n170));
BUF_X4 drc_ipo_c84 (.Z (out[19]), .A (drc_ipo_n168));
BUF_X4 drc_ipo_c83 (.Z (out[18]), .A (drc_ipo_n166));
BUF_X4 drc_ipo_c82 (.Z (out[17]), .A (drc_ipo_n164));
BUF_X4 drc_ipo_c81 (.Z (out[16]), .A (drc_ipo_n162));
BUF_X4 drc_ipo_c80 (.Z (out[15]), .A (drc_ipo_n160));
BUF_X4 drc_ipo_c79 (.Z (out[14]), .A (drc_ipo_n158));
BUF_X4 drc_ipo_c78 (.Z (out[13]), .A (drc_ipo_n156));
BUF_X4 drc_ipo_c77 (.Z (out[12]), .A (drc_ipo_n154));
BUF_X4 drc_ipo_c76 (.Z (out[11]), .A (drc_ipo_n152));
BUF_X4 drc_ipo_c75 (.Z (out[10]), .A (drc_ipo_n150));
BUF_X4 drc_ipo_c74 (.Z (out[9]), .A (drc_ipo_n148));
BUF_X4 drc_ipo_c73 (.Z (out[8]), .A (drc_ipo_n146));
BUF_X4 drc_ipo_c72 (.Z (out[7]), .A (drc_ipo_n144));
BUF_X4 drc_ipo_c71 (.Z (out[6]), .A (drc_ipo_n142));
BUF_X4 drc_ipo_c70 (.Z (out[5]), .A (drc_ipo_n140));
BUF_X4 drc_ipo_c69 (.Z (out[4]), .A (drc_ipo_n138));
BUF_X4 drc_ipo_c68 (.Z (out[3]), .A (drc_ipo_n136));
BUF_X4 drc_ipo_c67 (.Z (out[2]), .A (drc_ipo_n134));
BUF_X4 drc_ipo_c66 (.Z (out[1]), .A (drc_ipo_n132));
BUF_X4 drc_ipo_c65 (.Z (out[0]), .A (drc_ipo_n130));
CLKBUF_X3 CTS_L3_c99 (.Z (CTS_n194), .A (CTS_n195));

endmodule //registerNbits__2_5

module registerNbits__2_2 (clk_CTSPP_0, clk, reset, en, inp, out);

output [31:0] out;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTSPP_0;
wire drc_ipo_n192;
wire drc_ipo_n190;
wire drc_ipo_n188;
wire drc_ipo_n186;
wire drc_ipo_n184;
wire drc_ipo_n182;
wire drc_ipo_n180;
wire drc_ipo_n178;
wire drc_ipo_n176;
wire drc_ipo_n174;
wire drc_ipo_n172;
wire drc_ipo_n170;
wire drc_ipo_n168;
wire drc_ipo_n166;
wire drc_ipo_n164;
wire drc_ipo_n162;
wire drc_ipo_n160;
wire drc_ipo_n158;
wire drc_ipo_n156;
wire drc_ipo_n154;
wire drc_ipo_n152;
wire drc_ipo_n150;
wire drc_ipo_n148;
wire drc_ipo_n146;
wire drc_ipo_n144;
wire drc_ipo_n142;
wire drc_ipo_n140;
wire drc_ipo_n138;
wire drc_ipo_n136;
wire drc_ipo_n134;
wire drc_ipo_n132;
wire drc_ipo_n130;
wire n_0_0;
wire n_1;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n198;
wire CTS_n199;
wire CTS_n200;


AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (drc_ipo_n130), .CK (CTS_n200), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (drc_ipo_n132), .CK (CTS_n200), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (drc_ipo_n134), .CK (CTS_n200), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (drc_ipo_n136), .CK (CTS_n200), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (drc_ipo_n138), .CK (CTS_n200), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (drc_ipo_n140), .CK (CTS_n200), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (drc_ipo_n142), .CK (CTS_n200), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (drc_ipo_n144), .CK (CTS_n200), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (drc_ipo_n146), .CK (CTS_n199), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (drc_ipo_n148), .CK (CTS_n199), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (drc_ipo_n150), .CK (CTS_n199), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (drc_ipo_n152), .CK (CTS_n199), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (drc_ipo_n154), .CK (CTS_n199), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (drc_ipo_n156), .CK (CTS_n199), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (drc_ipo_n158), .CK (CTS_n199), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (drc_ipo_n160), .CK (CTS_n199), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (drc_ipo_n162), .CK (CTS_n199), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (drc_ipo_n164), .CK (CTS_n199), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (drc_ipo_n166), .CK (CTS_n200), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (drc_ipo_n168), .CK (CTS_n200), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (drc_ipo_n170), .CK (CTS_n200), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (drc_ipo_n172), .CK (CTS_n200), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (drc_ipo_n174), .CK (CTS_n200), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (drc_ipo_n176), .CK (CTS_n200), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (drc_ipo_n178), .CK (CTS_n200), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (drc_ipo_n180), .CK (CTS_n200), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (drc_ipo_n182), .CK (CTS_n200), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (drc_ipo_n184), .CK (CTS_n200), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (drc_ipo_n186), .CK (CTS_n200), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (drc_ipo_n188), .CK (CTS_n200), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (drc_ipo_n190), .CK (CTS_n200), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n192), .CK (CTS_n200), .D (n_33));
CLKGATETST_X4 clk_gate_out_reg (.GCK (CTS_n198), .CK (clk_CTSPP_0), .E (n_1), .SE (1'b0 ));
BUF_X4 drc_ipo_c96 (.Z (out[31]), .A (drc_ipo_n192));
BUF_X4 drc_ipo_c95 (.Z (out[30]), .A (drc_ipo_n190));
BUF_X4 drc_ipo_c94 (.Z (out[29]), .A (drc_ipo_n188));
BUF_X4 drc_ipo_c93 (.Z (out[28]), .A (drc_ipo_n186));
BUF_X4 drc_ipo_c92 (.Z (out[27]), .A (drc_ipo_n184));
BUF_X4 drc_ipo_c91 (.Z (out[26]), .A (drc_ipo_n182));
BUF_X4 drc_ipo_c90 (.Z (out[25]), .A (drc_ipo_n180));
BUF_X4 drc_ipo_c89 (.Z (out[24]), .A (drc_ipo_n178));
BUF_X4 drc_ipo_c88 (.Z (out[23]), .A (drc_ipo_n176));
BUF_X4 drc_ipo_c87 (.Z (out[22]), .A (drc_ipo_n174));
BUF_X4 drc_ipo_c86 (.Z (out[21]), .A (drc_ipo_n172));
BUF_X4 drc_ipo_c85 (.Z (out[20]), .A (drc_ipo_n170));
BUF_X4 drc_ipo_c84 (.Z (out[19]), .A (drc_ipo_n168));
BUF_X4 drc_ipo_c83 (.Z (out[18]), .A (drc_ipo_n166));
BUF_X4 drc_ipo_c82 (.Z (out[17]), .A (drc_ipo_n164));
BUF_X4 drc_ipo_c81 (.Z (out[16]), .A (drc_ipo_n162));
BUF_X4 drc_ipo_c80 (.Z (out[15]), .A (drc_ipo_n160));
BUF_X4 drc_ipo_c79 (.Z (out[14]), .A (drc_ipo_n158));
BUF_X4 drc_ipo_c78 (.Z (out[13]), .A (drc_ipo_n156));
BUF_X4 drc_ipo_c77 (.Z (out[12]), .A (drc_ipo_n154));
BUF_X4 drc_ipo_c76 (.Z (out[11]), .A (drc_ipo_n152));
BUF_X4 drc_ipo_c75 (.Z (out[10]), .A (drc_ipo_n150));
CLKBUF_X2 drc_ipo_c74 (.Z (out[9]), .A (drc_ipo_n148));
BUF_X4 drc_ipo_c73 (.Z (out[8]), .A (drc_ipo_n146));
BUF_X4 drc_ipo_c72 (.Z (out[7]), .A (drc_ipo_n144));
BUF_X4 drc_ipo_c71 (.Z (out[6]), .A (drc_ipo_n142));
BUF_X4 drc_ipo_c70 (.Z (out[5]), .A (drc_ipo_n140));
BUF_X4 drc_ipo_c69 (.Z (out[4]), .A (drc_ipo_n138));
BUF_X4 drc_ipo_c68 (.Z (out[3]), .A (drc_ipo_n136));
BUF_X4 drc_ipo_c67 (.Z (out[2]), .A (drc_ipo_n134));
BUF_X4 drc_ipo_c66 (.Z (out[1]), .A (drc_ipo_n132));
CLKBUF_X2 drc_ipo_c65 (.Z (out[0]), .A (drc_ipo_n130));
CLKBUF_X3 CTS_L3_c101 (.Z (CTS_n199), .A (CTS_n198));
CLKBUF_X3 CTS_L3_c102 (.Z (CTS_n200), .A (CTS_n198));

endmodule //registerNbits__2_2

module datapath (inputB, inputA, result);

output [63:0] result;
input [31:0] inputA;
input [31:0] inputB;
wire n_1030;
wire n_1045;
wire n_1053;
wire n_1052;
wire n_1040;
wire n_1046;
wire n_1069;
wire n_1068;
wire n_1056;
wire n_1074;
wire n_1073;
wire n_1084;
wire n_1077;
wire n_1098;
wire n_1097;
wire n_1072;
wire n_1103;
wire n_1102;
wire n_1078;
wire n_1092;
wire n_1127;
wire n_1126;
wire n_1113;
wire n_1106;
wire n_1132;
wire n_1131;
wire n_1128;
wire n_1101;
wire n_1137;
wire n_1136;
wire n_1114;
wire n_1107;
wire n_1160;
wire n_1159;
wire n_1154;
wire n_1147;
wire n_1165;
wire n_1164;
wire n_1161;
wire n_1130;
wire n_1170;
wire n_1169;
wire n_1135;
wire n_1166;
wire n_1175;
wire n_1174;
wire n_1141;
wire n_1192;
wire n_1206;
wire n_1205;
wire n_1178;
wire n_1163;
wire n_1211;
wire n_1210;
wire n_1168;
wire n_1207;
wire n_1216;
wire n_1215;
wire n_1173;
wire n_1221;
wire n_1220;
wire n_1186;
wire n_1179;
wire n_1252;
wire n_1251;
wire n_1244;
wire n_1238;
wire n_1257;
wire n_1256;
wire n_1224;
wire n_1253;
wire n_1262;
wire n_1261;
wire n_1214;
wire n_1258;
wire n_1267;
wire n_1266;
wire n_1219;
wire n_1272;
wire n_1271;
wire n_1239;
wire n_1232;
wire n_1302;
wire n_1301;
wire n_1245;
wire n_1296;
wire n_1307;
wire n_1306;
wire n_1282;
wire n_1275;
wire n_1312;
wire n_1311;
wire n_1303;
wire n_1260;
wire n_1317;
wire n_1316;
wire n_1313;
wire n_1308;
wire n_1322;
wire n_1321;
wire n_1270;
wire n_1327;
wire n_1326;
wire n_1283;
wire n_1276;
wire n_1365;
wire n_1364;
wire n_1351;
wire n_1344;
wire n_1370;
wire n_1369;
wire n_1330;
wire n_1366;
wire n_1375;
wire n_1374;
wire n_1310;
wire n_1315;
wire n_1380;
wire n_1379;
wire n_1320;
wire n_1376;
wire n_1385;
wire n_1384;
wire n_1325;
wire n_1390;
wire n_1389;
wire n_1345;
wire n_1338;
wire n_1428;
wire n_1427;
wire n_1359;
wire n_1420;
wire n_1433;
wire n_1432;
wire n_1407;
wire n_1400;
wire n_1438;
wire n_1437;
wire n_1368;
wire n_1429;
wire n_1443;
wire n_1442;
wire n_1378;
wire n_1439;
wire n_1448;
wire n_1447;
wire n_1444;
wire n_1383;
wire n_1453;
wire n_1452;
wire n_1449;
wire n_1458;
wire n_1457;
wire n_1415;
wire n_1408;
wire n_1495;
wire n_1494;
wire n_1394;
wire n_1431;
wire n_1500;
wire n_1499;
wire n_1489;
wire n_1482;
wire n_1505;
wire n_1504;
wire n_1468;
wire n_1461;
wire n_1510;
wire n_1509;
wire n_1441;
wire n_1436;
wire n_1515;
wire n_1514;
wire n_1446;
wire n_1511;
wire n_1520;
wire n_1519;
wire n_1516;
wire n_1451;
wire n_1525;
wire n_1524;
wire n_1456;
wire n_1530;
wire n_1529;
wire n_1476;
wire n_1469;
wire n_1575;
wire n_1574;
wire n_1498;
wire n_1561;
wire n_1580;
wire n_1579;
wire n_1547;
wire n_1540;
wire n_1585;
wire n_1584;
wire n_1503;
wire n_1576;
wire n_1590;
wire n_1589;
wire n_1508;
wire n_1513;
wire n_1595;
wire n_1594;
wire n_1581;
wire n_1518;
wire n_1600;
wire n_1599;
wire n_1523;
wire n_1596;
wire n_1605;
wire n_1604;
wire n_1528;
wire n_1610;
wire n_1609;
wire n_1555;
wire n_1548;
wire n_1655;
wire n_1654;
wire n_1534;
wire n_1578;
wire n_1660;
wire n_1659;
wire n_1647;
wire n_1641;
wire n_1665;
wire n_1664;
wire n_1627;
wire n_1620;
wire n_1670;
wire n_1669;
wire n_1656;
wire n_1588;
wire n_1675;
wire n_1674;
wire n_1661;
wire n_1593;
wire n_1680;
wire n_1679;
wire n_1666;
wire n_1676;
wire n_1685;
wire n_1684;
wire n_1681;
wire n_1603;
wire n_1690;
wire n_1689;
wire n_1608;
wire n_1695;
wire n_1694;
wire n_1642;
wire n_1635;
wire n_1739;
wire n_1738;
wire n_1621;
wire n_1614;
wire n_1744;
wire n_1743;
wire n_1648;
wire n_1733;
wire n_1749;
wire n_1748;
wire n_1719;
wire n_1712;
wire n_1754;
wire n_1753;
wire n_1698;
wire n_1663;
wire n_1759;
wire n_1758;
wire n_1740;
wire n_1673;
wire n_1764;
wire n_1763;
wire n_1678;
wire n_1755;
wire n_1769;
wire n_1768;
wire n_1760;
wire n_1765;
wire n_1774;
wire n_1773;
wire n_1688;
wire n_1770;
wire n_1779;
wire n_1778;
wire n_1693;
wire n_1784;
wire n_1783;
wire n_1720;
wire n_1713;
wire n_1836;
wire n_1835;
wire n_1699;
wire n_1742;
wire n_1841;
wire n_1840;
wire n_1815;
wire n_1808;
wire n_1846;
wire n_1845;
wire n_1794;
wire n_1787;
wire n_1851;
wire n_1850;
wire n_1837;
wire n_1829;
wire n_1856;
wire n_1855;
wire n_1752;
wire n_1842;
wire n_1861;
wire n_1860;
wire n_1762;
wire n_1852;
wire n_1866;
wire n_1865;
wire n_1857;
wire n_1772;
wire n_1871;
wire n_1870;
wire n_1777;
wire n_1867;
wire n_1876;
wire n_1875;
wire n_1782;
wire n_1877;
wire n_1881;
wire n_1880;
wire n_1816;
wire n_1809;
wire n_1933;
wire n_1932;
wire n_1795;
wire n_1788;
wire n_1938;
wire n_1937;
wire n_1830;
wire n_1925;
wire n_1943;
wire n_1942;
wire n_1912;
wire n_1905;
wire n_1948;
wire n_1947;
wire n_1891;
wire n_1884;
wire n_1953;
wire n_1952;
wire n_1934;
wire n_1849;
wire n_1958;
wire n_1957;
wire n_1854;
wire n_1859;
wire n_1963;
wire n_1962;
wire n_1949;
wire n_1944;
wire n_1968;
wire n_1967;
wire n_1959;
wire n_1869;
wire n_1973;
wire n_1972;
wire n_1969;
wire n_1874;
wire n_1978;
wire n_1977;
wire n_1879;
wire n_1979;
wire n_1983;
wire n_1982;
wire n_1920;
wire n_1913;
wire n_2034;
wire n_2033;
wire n_1899;
wire n_1892;
wire n_2039;
wire n_2038;
wire n_1936;
wire n_1926;
wire n_2044;
wire n_2043;
wire n_2021;
wire n_2014;
wire n_2049;
wire n_2048;
wire n_2000;
wire n_1993;
wire n_2054;
wire n_2053;
wire n_1941;
wire n_2040;
wire n_2059;
wire n_2058;
wire n_1951;
wire n_1946;
wire n_2064;
wire n_2063;
wire n_1961;
wire n_1956;
wire n_2069;
wire n_2068;
wire n_2050;
wire n_2065;
wire n_2074;
wire n_2073;
wire n_1966;
wire n_1971;
wire n_2079;
wire n_2078;
wire n_1976;
wire n_2075;
wire n_2084;
wire n_2083;
wire n_1981;
wire n_2089;
wire n_2088;
wire n_2015;
wire n_2008;
wire n_2148;
wire n_2147;
wire n_1994;
wire n_1987;
wire n_2153;
wire n_2152;
wire n_2037;
wire n_2134;
wire n_2158;
wire n_2157;
wire n_2120;
wire n_2113;
wire n_2163;
wire n_2162;
wire n_2099;
wire n_2092;
wire n_2168;
wire n_2167;
wire n_2149;
wire n_2141;
wire n_2173;
wire n_2172;
wire n_2052;
wire n_2047;
wire n_2178;
wire n_2177;
wire n_2169;
wire n_2164;
wire n_2183;
wire n_2182;
wire n_2067;
wire n_2179;
wire n_2188;
wire n_2187;
wire n_2072;
wire n_2077;
wire n_2193;
wire n_2192;
wire n_2082;
wire n_2189;
wire n_2198;
wire n_2197;
wire n_2087;
wire n_2199;
wire n_2203;
wire n_2202;
wire n_2128;
wire n_2121;
wire n_2262;
wire n_2261;
wire n_2107;
wire n_2100;
wire n_2267;
wire n_2266;
wire n_2151;
wire n_2142;
wire n_2272;
wire n_2271;
wire n_2248;
wire n_2241;
wire n_2277;
wire n_2276;
wire n_2227;
wire n_2220;
wire n_2282;
wire n_2281;
wire n_2206;
wire n_2156;
wire n_2287;
wire n_2286;
wire n_2263;
wire n_2166;
wire n_2292;
wire n_2291;
wire n_2273;
wire n_2176;
wire n_2297;
wire n_2296;
wire n_2283;
wire n_2278;
wire n_2302;
wire n_2301;
wire n_2181;
wire n_2293;
wire n_2307;
wire n_2306;
wire n_2298;
wire n_2191;
wire n_2312;
wire n_2311;
wire n_2308;
wire n_2196;
wire n_2317;
wire n_2316;
wire n_2201;
wire n_2318;
wire n_2322;
wire n_2321;
wire n_2249;
wire n_2242;
wire n_2380;
wire n_2379;
wire n_2228;
wire n_2221;
wire n_2385;
wire n_2384;
wire n_2207;
wire n_2270;
wire n_2390;
wire n_2389;
wire n_2255;
wire n_2374;
wire n_2395;
wire n_2394;
wire n_2360;
wire n_2353;
wire n_2400;
wire n_2399;
wire n_2339;
wire n_2332;
wire n_2405;
wire n_2404;
wire n_2386;
wire n_2381;
wire n_2410;
wire n_2409;
wire n_2280;
wire n_2275;
wire n_2415;
wire n_2414;
wire n_2295;
wire n_2290;
wire n_2420;
wire n_2419;
wire n_2401;
wire n_2396;
wire n_2425;
wire n_2424;
wire n_2416;
wire n_2411;
wire n_2430;
wire n_2429;
wire n_2421;
wire n_2310;
wire n_2435;
wire n_2434;
wire n_2431;
wire n_2315;
wire n_2440;
wire n_2439;
wire n_2320;
wire n_2441;
wire n_2445;
wire n_2444;
wire n_2361;
wire n_2354;
wire n_2511;
wire n_2510;
wire n_2340;
wire n_2333;
wire n_2516;
wire n_2515;
wire n_2388;
wire n_2383;
wire n_2521;
wire n_2520;
wire n_2490;
wire n_2483;
wire n_2526;
wire n_2525;
wire n_2469;
wire n_2462;
wire n_2531;
wire n_2530;
wire n_2448;
wire n_2393;
wire n_2536;
wire n_2535;
wire n_2512;
wire n_2504;
wire n_2541;
wire n_2540;
wire n_2403;
wire n_2398;
wire n_2546;
wire n_2545;
wire n_2413;
wire n_2532;
wire n_2551;
wire n_2550;
wire n_2537;
wire n_2418;
wire n_2556;
wire n_2555;
wire n_2542;
wire n_2423;
wire n_2561;
wire n_2560;
wire n_2433;
wire n_2552;
wire n_2566;
wire n_2565;
wire n_2562;
wire n_2438;
wire n_2571;
wire n_2570;
wire n_2443;
wire n_2572;
wire n_2576;
wire n_2575;
wire n_2491;
wire n_2484;
wire n_2642;
wire n_2641;
wire n_2470;
wire n_2463;
wire n_2647;
wire n_2646;
wire n_2449;
wire n_2519;
wire n_2652;
wire n_2651;
wire n_2505;
wire n_2634;
wire n_2657;
wire n_2656;
wire n_2621;
wire n_2614;
wire n_2662;
wire n_2661;
wire n_2600;
wire n_2593;
wire n_2667;
wire n_2666;
wire n_2579;
wire n_2648;
wire n_2672;
wire n_2671;
wire n_2534;
wire n_2529;
wire n_2677;
wire n_2676;
wire n_2653;
wire n_2544;
wire n_2682;
wire n_2681;
wire n_2668;
wire n_2663;
wire n_2687;
wire n_2686;
wire n_2549;
wire n_2678;
wire n_2692;
wire n_2691;
wire n_2554;
wire n_2683;
wire n_2697;
wire n_2696;
wire n_2564;
wire n_2688;
wire n_2702;
wire n_2701;
wire n_2569;
wire n_2698;
wire n_2707;
wire n_2706;
wire n_2574;
wire n_2712;
wire n_2711;
wire n_2629;
wire n_2622;
wire n_2777;
wire n_2776;
wire n_2608;
wire n_2601;
wire n_2782;
wire n_2781;
wire n_2587;
wire n_2580;
wire n_2787;
wire n_2786;
wire n_2645;
wire n_2635;
wire n_2792;
wire n_2791;
wire n_2764;
wire n_2757;
wire n_2797;
wire n_2796;
wire n_2743;
wire n_2736;
wire n_2802;
wire n_2801;
wire n_2722;
wire n_2715;
wire n_2807;
wire n_2806;
wire n_2788;
wire n_2783;
wire n_2812;
wire n_2811;
wire n_2670;
wire n_2665;
wire n_2817;
wire n_2816;
wire n_2793;
wire n_2680;
wire n_2822;
wire n_2821;
wire n_2808;
wire n_2803;
wire n_2827;
wire n_2826;
wire n_2685;
wire n_2818;
wire n_2832;
wire n_2831;
wire n_2690;
wire n_2823;
wire n_2837;
wire n_2836;
wire n_2828;
wire n_2700;
wire n_2842;
wire n_2841;
wire n_2838;
wire n_2705;
wire n_2847;
wire n_2846;
wire n_2710;
wire n_2848;
wire n_2852;
wire n_2851;
wire n_2758;
wire n_2751;
wire n_2925;
wire n_2924;
wire n_2737;
wire n_2730;
wire n_2930;
wire n_2929;
wire n_2716;
wire n_2785;
wire n_2935;
wire n_2934;
wire n_2911;
wire n_2904;
wire n_2940;
wire n_2939;
wire n_2890;
wire n_2883;
wire n_2945;
wire n_2944;
wire n_2869;
wire n_2862;
wire n_2950;
wire n_2949;
wire n_2790;
wire n_2931;
wire n_2955;
wire n_2954;
wire n_2918;
wire n_2805;
wire n_2960;
wire n_2959;
wire n_2795;
wire n_2810;
wire n_2965;
wire n_2964;
wire n_2820;
wire n_2815;
wire n_2970;
wire n_2969;
wire n_2946;
wire n_2941;
wire n_2975;
wire n_2974;
wire n_2961;
wire n_2956;
wire n_2980;
wire n_2979;
wire n_2966;
wire n_2971;
wire n_2985;
wire n_2984;
wire n_2976;
wire n_2840;
wire n_2990;
wire n_2989;
wire n_2986;
wire n_2845;
wire n_2995;
wire n_2994;
wire n_2850;
wire n_2996;
wire n_3000;
wire n_2999;
wire n_2905;
wire n_2898;
wire n_3073;
wire n_3072;
wire n_2884;
wire n_2877;
wire n_3078;
wire n_3077;
wire n_2863;
wire n_2856;
wire n_3083;
wire n_3082;
wire n_2928;
wire n_2919;
wire n_3088;
wire n_3087;
wire n_3059;
wire n_3052;
wire n_3093;
wire n_3092;
wire n_3038;
wire n_3031;
wire n_3098;
wire n_3097;
wire n_3017;
wire n_3010;
wire n_3103;
wire n_3102;
wire n_2938;
wire n_3084;
wire n_3108;
wire n_3107;
wire n_3074;
wire n_2953;
wire n_3113;
wire n_3112;
wire n_2943;
wire n_3089;
wire n_3118;
wire n_3117;
wire n_2958;
wire n_3104;
wire n_3123;
wire n_3122;
wire n_3094;
wire n_2968;
wire n_3128;
wire n_3127;
wire n_3109;
wire n_2973;
wire n_3133;
wire n_3132;
wire n_3119;
wire n_2983;
wire n_3138;
wire n_3137;
wire n_3129;
wire n_2988;
wire n_3143;
wire n_3142;
wire n_3139;
wire n_2993;
wire n_3148;
wire n_3147;
wire n_2998;
wire n_3149;
wire n_3153;
wire n_3152;
wire n_3060;
wire n_3053;
wire n_3225;
wire n_3224;
wire n_3039;
wire n_3032;
wire n_3230;
wire n_3229;
wire n_3018;
wire n_3011;
wire n_3235;
wire n_3234;
wire n_3081;
wire n_3076;
wire n_3240;
wire n_3239;
wire n_3219;
wire n_3212;
wire n_3245;
wire n_3244;
wire n_3198;
wire n_3191;
wire n_3250;
wire n_3249;
wire n_3177;
wire n_3170;
wire n_3255;
wire n_3254;
wire n_3156;
wire n_3086;
wire n_3260;
wire n_3259;
wire n_3231;
wire n_3226;
wire n_3265;
wire n_3264;
wire n_3101;
wire n_3096;
wire n_3270;
wire n_3269;
wire n_3241;
wire n_3116;
wire n_3275;
wire n_3274;
wire n_3256;
wire n_3251;
wire n_3280;
wire n_3279;
wire n_3261;
wire n_3121;
wire n_3285;
wire n_3284;
wire n_3266;
wire n_3126;
wire n_3290;
wire n_3289;
wire n_3131;
wire n_3136;
wire n_3295;
wire n_3294;
wire n_3286;
wire n_3291;
wire n_3300;
wire n_3299;
wire n_3146;
wire n_3296;
wire n_3305;
wire n_3304;
wire n_3151;
wire n_3306;
wire n_3310;
wire n_3309;
wire n_3206;
wire n_3199;
wire n_3390;
wire n_3389;
wire n_3185;
wire n_3178;
wire n_3395;
wire n_3394;
wire n_3164;
wire n_3157;
wire n_3400;
wire n_3399;
wire n_3233;
wire n_3228;
wire n_3405;
wire n_3404;
wire n_3369;
wire n_3362;
wire n_3410;
wire n_3409;
wire n_3348;
wire n_3341;
wire n_3415;
wire n_3414;
wire n_3327;
wire n_3320;
wire n_3420;
wire n_3419;
wire n_3243;
wire n_3401;
wire n_3425;
wire n_3424;
wire n_3391;
wire n_3383;
wire n_3430;
wire n_3429;
wire n_3253;
wire n_3248;
wire n_3435;
wire n_3434;
wire n_3273;
wire n_3268;
wire n_3440;
wire n_3439;
wire n_3421;
wire n_3416;
wire n_3445;
wire n_3444;
wire n_3278;
wire n_3436;
wire n_3450;
wire n_3449;
wire n_3426;
wire n_3283;
wire n_3455;
wire n_3454;
wire n_3288;
wire n_3446;
wire n_3460;
wire n_3459;
wire n_3456;
wire n_3451;
wire n_3465;
wire n_3464;
wire n_3303;
wire n_3461;
wire n_3470;
wire n_3469;
wire n_3308;
wire n_3471;
wire n_3475;
wire n_3474;
wire n_3370;
wire n_3363;
wire n_3556;
wire n_3555;
wire n_3349;
wire n_3342;
wire n_3561;
wire n_3560;
wire n_3328;
wire n_3321;
wire n_3566;
wire n_3565;
wire n_3398;
wire n_3393;
wire n_3571;
wire n_3570;
wire n_3549;
wire n_3542;
wire n_3576;
wire n_3575;
wire n_3528;
wire n_3521;
wire n_3581;
wire n_3580;
wire n_3507;
wire n_3500;
wire n_3586;
wire n_3585;
wire n_3486;
wire n_3477;
wire n_3591;
wire n_3590;
wire n_3567;
wire n_3562;
wire n_3596;
wire n_3595;
wire n_3423;
wire n_3418;
wire n_3601;
wire n_3600;
wire n_3408;
wire n_3572;
wire n_3606;
wire n_3605;
wire n_3428;
wire n_3592;
wire n_3611;
wire n_3610;
wire n_3582;
wire n_3577;
wire n_3616;
wire n_3615;
wire n_3438;
wire n_3602;
wire n_3621;
wire n_3620;
wire n_3448;
wire n_3607;
wire n_3626;
wire n_3625;
wire n_3617;
wire n_3612;
wire n_3631;
wire n_3630;
wire n_3622;
wire n_3463;
wire n_3636;
wire n_3635;
wire n_3468;
wire n_3632;
wire n_3641;
wire n_3640;
wire n_3473;
wire n_3642;
wire n_3646;
wire n_3645;
wire n_3536;
wire n_3529;
wire n_3723;
wire n_3722;
wire n_3515;
wire n_3508;
wire n_3728;
wire n_3727;
wire n_3494;
wire n_3487;
wire n_3733;
wire n_3732;
wire n_3569;
wire n_3564;
wire n_3738;
wire n_3737;
wire n_3550;
wire n_3716;
wire n_3743;
wire n_3742;
wire n_3702;
wire n_3695;
wire n_3748;
wire n_3747;
wire n_3681;
wire n_3674;
wire n_3753;
wire n_3752;
wire n_3660;
wire n_3653;
wire n_3758;
wire n_3757;
wire n_3574;
wire n_3734;
wire n_3763;
wire n_3762;
wire n_3724;
wire n_3589;
wire n_3768;
wire n_3767;
wire n_3579;
wire n_3594;
wire n_3773;
wire n_3772;
wire n_3604;
wire n_3599;
wire n_3778;
wire n_3777;
wire n_3754;
wire n_3749;
wire n_3783;
wire n_3782;
wire n_3609;
wire n_3769;
wire n_3788;
wire n_3787;
wire n_3614;
wire n_3774;
wire n_3793;
wire n_3792;
wire n_3779;
wire n_3624;
wire n_3798;
wire n_3797;
wire n_3629;
wire n_3789;
wire n_3803;
wire n_3802;
wire n_3634;
wire n_3799;
wire n_3808;
wire n_3807;
wire n_3804;
wire n_3809;
wire n_3813;
wire n_3812;
wire n_3710;
wire n_3703;
wire n_3890;
wire n_3889;
wire n_3689;
wire n_3682;
wire n_3895;
wire n_3894;
wire n_3668;
wire n_3661;
wire n_3900;
wire n_3899;
wire n_3649;
wire n_3736;
wire n_3905;
wire n_3904;
wire n_3726;
wire n_3717;
wire n_3910;
wire n_3909;
wire n_3876;
wire n_3869;
wire n_3915;
wire n_3914;
wire n_3855;
wire n_3848;
wire n_3920;
wire n_3919;
wire n_3834;
wire n_3827;
wire n_3925;
wire n_3924;
wire n_3741;
wire n_3901;
wire n_3930;
wire n_3929;
wire n_3891;
wire n_3761;
wire n_3935;
wire n_3934;
wire n_3751;
wire n_3746;
wire n_3940;
wire n_3939;
wire n_3906;
wire n_3771;
wire n_3945;
wire n_3944;
wire n_3926;
wire n_3921;
wire n_3950;
wire n_3949;
wire n_3776;
wire n_3941;
wire n_3955;
wire n_3954;
wire n_3931;
wire n_3786;
wire n_3960;
wire n_3959;
wire n_3946;
wire n_3791;
wire n_3965;
wire n_3964;
wire n_3951;
wire n_3961;
wire n_3970;
wire n_3969;
wire n_3801;
wire n_3966;
wire n_3975;
wire n_3974;
wire n_3971;
wire n_3811;
wire n_3980;
wire n_3979;
wire n_3877;
wire n_3870;
wire n_4057;
wire n_4056;
wire n_3856;
wire n_3849;
wire n_4062;
wire n_4061;
wire n_3835;
wire n_3828;
wire n_4067;
wire n_4066;
wire n_3903;
wire n_3898;
wire n_4072;
wire n_4071;
wire n_4050;
wire n_4043;
wire n_4077;
wire n_4076;
wire n_4029;
wire n_4022;
wire n_4082;
wire n_4081;
wire n_4008;
wire n_4001;
wire n_4087;
wire n_4086;
wire n_3985;
wire n_3908;
wire n_4092;
wire n_4091;
wire n_4063;
wire n_4058;
wire n_4097;
wire n_4096;
wire n_3923;
wire n_3918;
wire n_4102;
wire n_4101;
wire n_4073;
wire n_3938;
wire n_4107;
wire n_4106;
wire n_4088;
wire n_4083;
wire n_4112;
wire n_4111;
wire n_4093;
wire n_3948;
wire n_4117;
wire n_4116;
wire n_4103;
wire n_4098;
wire n_4122;
wire n_4121;
wire n_4108;
wire n_3963;
wire n_4127;
wire n_4126;
wire n_4113;
wire n_4118;
wire n_4132;
wire n_4131;
wire n_4123;
wire n_4128;
wire n_4137;
wire n_4136;
wire n_4133;
wire n_3978;
wire n_4142;
wire n_4141;
wire n_384;
wire n_4044;
wire n_4211;
wire n_4210;
wire n_4030;
wire n_4023;
wire n_4216;
wire n_4215;
wire n_4009;
wire n_4002;
wire n_4221;
wire n_4220;
wire n_3986;
wire n_4070;
wire n_4226;
wire n_4225;
wire n_4060;
wire n_4051;
wire n_4231;
wire n_4230;
wire n_4198;
wire n_4191;
wire n_4236;
wire n_4235;
wire n_4177;
wire n_4170;
wire n_4241;
wire n_4240;
wire n_4156;
wire n_4147;
wire n_4246;
wire n_4245;
wire n_4222;
wire n_4217;
wire n_4251;
wire n_4250;
wire n_4090;
wire n_4085;
wire n_4256;
wire n_4255;
wire n_4232;
wire n_4227;
wire n_4261;
wire n_4260;
wire n_4100;
wire n_4095;
wire n_4266;
wire n_4265;
wire n_4242;
wire n_4237;
wire n_4271;
wire n_4270;
wire n_4257;
wire n_4252;
wire n_4276;
wire n_4275;
wire n_4120;
wire n_4267;
wire n_4281;
wire n_4280;
wire n_4125;
wire n_4272;
wire n_4286;
wire n_4285;
wire n_4277;
wire n_4135;
wire n_4291;
wire n_4290;
wire n_4287;
wire n_4140;
wire n_4296;
wire n_4295;
wire n_4206;
wire n_4199;
wire n_4366;
wire n_4365;
wire n_4185;
wire n_4178;
wire n_4371;
wire n_4370;
wire n_4164;
wire n_4157;
wire n_4376;
wire n_4375;
wire n_4224;
wire n_4219;
wire n_4381;
wire n_4380;
wire n_4358;
wire n_4352;
wire n_4386;
wire n_4385;
wire n_4338;
wire n_4331;
wire n_4391;
wire n_4390;
wire n_4317;
wire n_4310;
wire n_4396;
wire n_4395;
wire n_4229;
wire n_4377;
wire n_4401;
wire n_4400;
wire n_4367;
wire n_4244;
wire n_4406;
wire n_4405;
wire n_4234;
wire n_4249;
wire n_4411;
wire n_4410;
wire n_4259;
wire n_4254;
wire n_4416;
wire n_4415;
wire n_4392;
wire n_4387;
wire n_4421;
wire n_4420;
wire n_4407;
wire n_4402;
wire n_4426;
wire n_4425;
wire n_4412;
wire n_4274;
wire n_4431;
wire n_4430;
wire n_4279;
wire n_4422;
wire n_4436;
wire n_4435;
wire n_4427;
wire n_4432;
wire n_4441;
wire n_4440;
wire n_4437;
wire n_4294;
wire n_4446;
wire n_4445;
wire n_4353;
wire n_4346;
wire n_4516;
wire n_4515;
wire n_4332;
wire n_4325;
wire n_4521;
wire n_4520;
wire n_4311;
wire n_4302;
wire n_4526;
wire n_4525;
wire n_4374;
wire n_4369;
wire n_4531;
wire n_4530;
wire n_4502;
wire n_4495;
wire n_4536;
wire n_4535;
wire n_4481;
wire n_4474;
wire n_4541;
wire n_4540;
wire n_4460;
wire n_4451;
wire n_4546;
wire n_4545;
wire n_4527;
wire n_4522;
wire n_4551;
wire n_4550;
wire n_4399;
wire n_4394;
wire n_4556;
wire n_4555;
wire n_4532;
wire n_4409;
wire n_4561;
wire n_4560;
wire n_4547;
wire n_4542;
wire n_4566;
wire n_4565;
wire n_4414;
wire n_4557;
wire n_4571;
wire n_4570;
wire n_4419;
wire n_4424;
wire n_4576;
wire n_4575;
wire n_4429;
wire n_4567;
wire n_4581;
wire n_4580;
wire n_4572;
wire n_4577;
wire n_4586;
wire n_4585;
wire n_4444;
wire n_4582;
wire n_4591;
wire n_4590;
wire n_383;
wire n_4503;
wire n_4653;
wire n_4652;
wire n_4489;
wire n_4482;
wire n_4658;
wire n_4657;
wire n_4468;
wire n_4461;
wire n_4663;
wire n_4662;
wire n_4524;
wire n_4519;
wire n_4668;
wire n_4667;
wire n_4647;
wire n_4640;
wire n_4673;
wire n_4672;
wire n_4626;
wire n_4619;
wire n_4678;
wire n_4677;
wire n_4605;
wire n_4596;
wire n_4683;
wire n_4682;
wire n_4664;
wire n_4659;
wire n_4688;
wire n_4687;
wire n_4544;
wire n_4539;
wire n_4693;
wire n_4692;
wire n_4549;
wire n_4669;
wire n_4698;
wire n_4697;
wire n_4554;
wire n_4684;
wire n_4703;
wire n_4702;
wire n_4674;
wire n_4564;
wire n_4708;
wire n_4707;
wire n_4689;
wire n_4569;
wire n_4713;
wire n_4712;
wire n_4574;
wire n_4704;
wire n_4718;
wire n_4717;
wire n_4579;
wire n_4714;
wire n_4723;
wire n_4722;
wire n_4589;
wire n_4719;
wire n_4728;
wire n_4727;
wire n_4648;
wire n_4641;
wire n_4791;
wire n_4790;
wire n_4627;
wire n_4620;
wire n_4796;
wire n_4795;
wire n_4606;
wire n_4597;
wire n_4801;
wire n_4800;
wire n_4661;
wire n_4656;
wire n_4806;
wire n_4805;
wire n_4777;
wire n_4770;
wire n_4811;
wire n_4810;
wire n_4756;
wire n_4749;
wire n_4816;
wire n_4815;
wire n_4733;
wire n_4671;
wire n_4821;
wire n_4820;
wire n_4797;
wire n_4792;
wire n_4826;
wire n_4825;
wire n_4676;
wire n_4686;
wire n_4831;
wire n_4830;
wire n_4696;
wire n_4691;
wire n_4836;
wire n_4835;
wire n_4812;
wire n_4822;
wire n_4841;
wire n_4840;
wire n_4827;
wire n_4706;
wire n_4846;
wire n_4845;
wire n_4837;
wire n_4711;
wire n_4851;
wire n_4850;
wire n_4716;
wire n_4847;
wire n_4856;
wire n_4855;
wire n_4852;
wire n_4726;
wire n_4861;
wire n_4860;
wire n_4778;
wire n_4771;
wire n_4924;
wire n_4923;
wire n_4757;
wire n_4750;
wire n_4929;
wire n_4928;
wire n_4734;
wire n_4799;
wire n_4934;
wire n_4933;
wire n_4917;
wire n_4910;
wire n_4939;
wire n_4938;
wire n_4896;
wire n_4889;
wire n_4944;
wire n_4943;
wire n_4875;
wire n_4866;
wire n_4949;
wire n_4948;
wire n_4930;
wire n_4925;
wire n_4954;
wire n_4953;
wire n_4814;
wire n_4809;
wire n_4959;
wire n_4958;
wire n_4829;
wire n_4824;
wire n_4964;
wire n_4963;
wire n_4945;
wire n_4940;
wire n_4969;
wire n_4968;
wire n_4960;
wire n_4955;
wire n_4974;
wire n_4973;
wire n_4844;
wire n_4965;
wire n_4979;
wire n_4978;
wire n_4970;
wire n_4975;
wire n_4984;
wire n_4983;
wire n_4980;
wire n_4859;
wire n_4989;
wire n_4988;
wire n_382;
wire n_4911;
wire n_5044;
wire n_5043;
wire n_4897;
wire n_4890;
wire n_5049;
wire n_5048;
wire n_4876;
wire n_4867;
wire n_5054;
wire n_5053;
wire n_4927;
wire n_4918;
wire n_5059;
wire n_5058;
wire n_5031;
wire n_5024;
wire n_5064;
wire n_5063;
wire n_5010;
wire n_5003;
wire n_5069;
wire n_5068;
wire n_4937;
wire n_5055;
wire n_5074;
wire n_5073;
wire n_5045;
wire n_4947;
wire n_5079;
wire n_5078;
wire n_4952;
wire n_5060;
wire n_5084;
wire n_5083;
wire n_5070;
wire n_5065;
wire n_5089;
wire n_5088;
wire n_5080;
wire n_5075;
wire n_5094;
wire n_5093;
wire n_4972;
wire n_5085;
wire n_5099;
wire n_5098;
wire n_5090;
wire n_4982;
wire n_5104;
wire n_5103;
wire n_5100;
wire n_4987;
wire n_5109;
wire n_5108;
wire n_5039;
wire n_5032;
wire n_5165;
wire n_5164;
wire n_5018;
wire n_5011;
wire n_5170;
wire n_5169;
wire n_4995;
wire n_5052;
wire n_5175;
wire n_5174;
wire n_5157;
wire n_5151;
wire n_5180;
wire n_5179;
wire n_5137;
wire n_5130;
wire n_5185;
wire n_5184;
wire n_5114;
wire n_5057;
wire n_5190;
wire n_5189;
wire n_5166;
wire n_5072;
wire n_5195;
wire n_5194;
wire n_5062;
wire n_5176;
wire n_5200;
wire n_5199;
wire n_5077;
wire n_5186;
wire n_5205;
wire n_5204;
wire n_5191;
wire n_5087;
wire n_5210;
wire n_5209;
wire n_5092;
wire n_5201;
wire n_5215;
wire n_5214;
wire n_5206;
wire n_5211;
wire n_5220;
wire n_5219;
wire n_5216;
wire n_5107;
wire n_5225;
wire n_5224;
wire n_5152;
wire n_5145;
wire n_5281;
wire n_5280;
wire n_5131;
wire n_5124;
wire n_5286;
wire n_5285;
wire n_5173;
wire n_5168;
wire n_5291;
wire n_5290;
wire n_5267;
wire n_5260;
wire n_5296;
wire n_5295;
wire n_5246;
wire n_5239;
wire n_5301;
wire n_5300;
wire n_5178;
wire n_5287;
wire n_5306;
wire n_5305;
wire n_5188;
wire n_5183;
wire n_5311;
wire n_5310;
wire n_5198;
wire n_5193;
wire n_5316;
wire n_5315;
wire n_5297;
wire n_5203;
wire n_5321;
wire n_5320;
wire n_5307;
wire n_5208;
wire n_5326;
wire n_5325;
wire n_5213;
wire n_5322;
wire n_5331;
wire n_5330;
wire n_5327;
wire n_5223;
wire n_5336;
wire n_5335;
wire n_447;
wire n_5268;
wire n_5384;
wire n_5383;
wire n_5254;
wire n_5247;
wire n_5389;
wire n_5388;
wire n_5231;
wire n_5289;
wire n_5394;
wire n_5393;
wire n_5275;
wire n_5378;
wire n_5399;
wire n_5398;
wire n_5364;
wire n_5357;
wire n_5404;
wire n_5403;
wire n_5341;
wire n_5390;
wire n_5409;
wire n_5408;
wire n_5304;
wire n_5299;
wire n_5414;
wire n_5413;
wire n_5395;
wire n_5309;
wire n_5419;
wire n_5418;
wire n_5400;
wire n_5314;
wire n_5424;
wire n_5423;
wire n_5410;
wire n_5319;
wire n_5429;
wire n_5428;
wire n_5324;
wire n_5425;
wire n_5434;
wire n_5433;
wire n_5430;
wire n_5334;
wire n_5439;
wire n_5438;
wire n_5379;
wire n_5372;
wire n_5488;
wire n_5487;
wire n_5358;
wire n_5351;
wire n_5493;
wire n_5492;
wire n_5392;
wire n_5387;
wire n_5498;
wire n_5497;
wire n_5474;
wire n_5467;
wire n_5503;
wire n_5502;
wire n_5453;
wire n_5444;
wire n_5508;
wire n_5507;
wire n_5494;
wire n_5489;
wire n_5513;
wire n_5512;
wire n_5402;
wire n_5499;
wire n_5518;
wire n_5517;
wire n_5412;
wire n_5509;
wire n_5523;
wire n_5522;
wire n_5514;
wire n_5422;
wire n_5528;
wire n_5527;
wire n_5427;
wire n_5524;
wire n_5533;
wire n_5532;
wire n_5529;
wire n_5437;
wire n_5538;
wire n_5537;
wire n_5475;
wire n_5468;
wire n_5587;
wire n_5586;
wire n_5454;
wire n_5445;
wire n_5592;
wire n_5591;
wire n_5491;
wire n_5580;
wire n_5597;
wire n_5596;
wire n_5566;
wire n_5559;
wire n_5602;
wire n_5601;
wire n_5543;
wire n_5593;
wire n_5607;
wire n_5606;
wire n_5506;
wire n_5501;
wire n_5612;
wire n_5611;
wire n_5516;
wire n_5603;
wire n_5617;
wire n_5616;
wire n_5521;
wire n_5613;
wire n_5622;
wire n_5621;
wire n_5526;
wire n_5618;
wire n_5627;
wire n_5626;
wire n_5623;
wire n_5536;
wire n_5632;
wire n_5631;
wire n_543;
wire n_5574;
wire n_5673;
wire n_5672;
wire n_5560;
wire n_5553;
wire n_5678;
wire n_5677;
wire n_5590;
wire n_5581;
wire n_5683;
wire n_5682;
wire n_5660;
wire n_5653;
wire n_5688;
wire n_5687;
wire n_5637;
wire n_5595;
wire n_5693;
wire n_5692;
wire n_5674;
wire n_5605;
wire n_5698;
wire n_5697;
wire n_5684;
wire n_5610;
wire n_5703;
wire n_5702;
wire n_5689;
wire n_5694;
wire n_5708;
wire n_5707;
wire n_5620;
wire n_5704;
wire n_5713;
wire n_5712;
wire n_5709;
wire n_5630;
wire n_5718;
wire n_5717;
wire n_5668;
wire n_5661;
wire n_5760;
wire n_5759;
wire n_5647;
wire n_5638;
wire n_5765;
wire n_5764;
wire n_5676;
wire n_5752;
wire n_1;
wire n_0;
wire n_5739;
wire n_5732;
wire n_3;
wire n_2;
wire n_5766;
wire n_5761;
wire n_5;
wire n_4;
wire n_5686;
wire n_5701;
wire n_7;
wire n_6;
wire n_381;
wire n_380;
wire n_9;
wire n_8;
wire n_379;
wire n_378;
wire n_11;
wire n_10;
wire n_377;
wire n_5716;
wire n_13;
wire n_12;
wire n_5747;
wire n_5740;
wire n_15;
wire n_14;
wire n_5724;
wire n_5763;
wire n_17;
wire n_16;
wire n_376;
wire n_375;
wire n_19;
wire n_18;
wire n_374;
wire n_373;
wire n_21;
wire n_20;
wire n_372;
wire n_371;
wire n_23;
wire n_22;
wire n_370;
wire n_369;
wire n_25;
wire n_24;
wire n_368;
wire n_367;
wire n_27;
wire n_26;
wire n_366;
wire n_365;
wire n_29;
wire n_28;
wire n_639;
wire n_364;
wire n_31;
wire n_30;
wire n_363;
wire n_362;
wire n_33;
wire n_32;
wire n_361;
wire n_360;
wire n_35;
wire n_34;
wire n_359;
wire n_358;
wire n_37;
wire n_36;
wire n_357;
wire n_356;
wire n_39;
wire n_38;
wire n_355;
wire n_354;
wire n_41;
wire n_40;
wire n_353;
wire n_352;
wire n_43;
wire n_42;
wire n_351;
wire n_350;
wire n_45;
wire n_44;
wire n_349;
wire n_348;
wire n_47;
wire n_46;
wire n_347;
wire n_346;
wire n_49;
wire n_48;
wire n_345;
wire n_344;
wire n_51;
wire n_50;
wire n_343;
wire n_342;
wire n_53;
wire n_52;
wire n_341;
wire n_340;
wire n_55;
wire n_54;
wire n_339;
wire n_338;
wire n_57;
wire n_56;
wire n_337;
wire n_336;
wire n_59;
wire n_58;
wire n_335;
wire n_334;
wire n_61;
wire n_60;
wire n_333;
wire n_332;
wire n_63;
wire n_62;
wire n_331;
wire n_330;
wire n_65;
wire n_64;
wire n_329;
wire n_328;
wire n_67;
wire n_66;
wire n_327;
wire n_326;
wire n_69;
wire n_68;
wire n_325;
wire n_324;
wire n_71;
wire n_70;
wire n_735;
wire n_323;
wire n_73;
wire n_72;
wire n_322;
wire n_321;
wire n_75;
wire n_74;
wire n_320;
wire n_319;
wire n_77;
wire n_76;
wire n_318;
wire n_317;
wire n_79;
wire n_78;
wire n_316;
wire n_315;
wire n_81;
wire n_80;
wire n_314;
wire n_313;
wire n_83;
wire n_82;
wire n_312;
wire n_311;
wire n_85;
wire n_84;
wire n_310;
wire n_309;
wire n_87;
wire n_86;
wire n_308;
wire n_307;
wire n_89;
wire n_88;
wire n_306;
wire n_305;
wire n_91;
wire n_90;
wire n_304;
wire n_303;
wire n_93;
wire n_92;
wire n_302;
wire n_301;
wire n_95;
wire n_94;
wire n_300;
wire n_299;
wire n_97;
wire n_96;
wire n_298;
wire n_297;
wire n_99;
wire n_98;
wire n_296;
wire n_295;
wire n_101;
wire n_100;
wire n_831;
wire n_294;
wire n_103;
wire n_102;
wire n_293;
wire n_292;
wire n_105;
wire n_104;
wire n_291;
wire n_290;
wire n_107;
wire n_106;
wire n_289;
wire n_288;
wire n_109;
wire n_108;
wire n_287;
wire n_286;
wire n_111;
wire n_110;
wire n_285;
wire n_284;
wire n_113;
wire n_112;
wire n_283;
wire n_282;
wire n_115;
wire n_114;
wire n_281;
wire n_280;
wire n_117;
wire n_116;
wire n_279;
wire n_278;
wire n_119;
wire n_118;
wire n_927;
wire n_277;
wire n_121;
wire n_120;
wire n_276;
wire n_275;
wire n_123;
wire n_122;
wire n_274;
wire n_273;
wire n_125;
wire n_124;
wire n_1022;
wire n_991;
wire n_127;
wire n_126;
wire n_1034;
wire n_1029;
wire n_129;
wire n_128;
wire n_1039;
wire n_131;
wire n_130;
wire n_1070;
wire n_133;
wire n_132;
wire n_1099;
wire n_135;
wire n_134;
wire n_1133;
wire n_137;
wire n_136;
wire n_1171;
wire n_139;
wire n_138;
wire n_1217;
wire n_141;
wire n_140;
wire n_1268;
wire n_143;
wire n_142;
wire n_1323;
wire n_145;
wire n_144;
wire n_1386;
wire n_147;
wire n_146;
wire n_1454;
wire n_149;
wire n_148;
wire n_1526;
wire n_151;
wire n_150;
wire n_1606;
wire n_153;
wire n_152;
wire n_1691;
wire n_155;
wire n_154;
wire n_1780;
wire n_157;
wire n_156;
wire n_159;
wire n_158;
wire n_161;
wire n_160;
wire n_2085;
wire n_163;
wire n_162;
wire n_165;
wire n_164;
wire n_167;
wire n_166;
wire n_169;
wire n_168;
wire n_171;
wire n_170;
wire n_2708;
wire n_173;
wire n_172;
wire n_175;
wire n_174;
wire n_177;
wire n_176;
wire n_179;
wire n_178;
wire n_181;
wire n_180;
wire n_183;
wire n_182;
wire n_185;
wire n_184;
wire n_3814;
wire n_187;
wire n_186;
wire n_3816;
wire n_3981;
wire n_189;
wire n_188;
wire n_3983;
wire n_4143;
wire n_191;
wire n_190;
wire n_4297;
wire n_4145;
wire n_193;
wire n_192;
wire n_4299;
wire n_4447;
wire n_195;
wire n_194;
wire n_4449;
wire n_4592;
wire n_197;
wire n_196;
wire n_4594;
wire n_4729;
wire n_199;
wire n_198;
wire n_4731;
wire n_4862;
wire n_201;
wire n_200;
wire n_4864;
wire n_4990;
wire n_203;
wire n_202;
wire n_4992;
wire n_5110;
wire n_205;
wire n_204;
wire n_5112;
wire n_5226;
wire n_207;
wire n_206;
wire n_5228;
wire n_5337;
wire n_209;
wire n_208;
wire n_5339;
wire n_5440;
wire n_211;
wire n_210;
wire n_5442;
wire n_5539;
wire n_213;
wire n_212;
wire n_5541;
wire n_5633;
wire n_215;
wire n_214;
wire n_5635;
wire n_5719;
wire n_217;
wire n_216;
wire n_5721;
wire n_272;
wire n_219;
wire n_218;
wire n_271;
wire n_270;
wire n_221;
wire n_220;
wire n_269;
wire n_268;
wire n_223;
wire n_222;
wire n_267;
wire n_266;
wire n_225;
wire n_224;
wire n_265;
wire n_264;
wire n_227;
wire n_226;
wire n_263;
wire n_262;
wire n_229;
wire n_228;
wire n_261;
wire n_260;
wire n_231;
wire n_230;
wire n_259;
wire n_258;
wire n_233;
wire n_232;
wire n_257;
wire n_256;
wire n_235;
wire n_234;
wire n_255;
wire n_254;
wire n_237;
wire n_236;
wire n_253;
wire n_252;
wire n_239;
wire n_238;
wire n_251;
wire n_250;
wire n_241;
wire n_240;
wire n_249;
wire n_248;
wire n_243;
wire n_242;
wire n_247;
wire n_246;
wire n_245;
wire n_244;
wire n_385;
wire n_386;
wire n_5742;
wire n_387;
wire n_454;
wire n_388;
wire n_390;
wire n_389;
wire n_392;
wire n_391;
wire n_393;
wire n_460;
wire n_394;
wire n_461;
wire n_484;
wire n_462;
wire n_395;
wire n_397;
wire n_396;
wire n_398;
wire n_465;
wire n_476;
wire n_399;
wire n_401;
wire n_400;
wire n_403;
wire n_402;
wire n_404;
wire n_508;
wire n_405;
wire n_406;
wire n_535;
wire n_407;
wire n_409;
wire n_408;
wire n_410;
wire n_561;
wire n_590;
wire n_411;
wire n_412;
wire n_624;
wire n_413;
wire n_415;
wire n_414;
wire n_416;
wire n_671;
wire n_700;
wire n_417;
wire n_418;
wire n_748;
wire n_419;
wire n_420;
wire n_793;
wire n_421;
wire n_422;
wire n_840;
wire n_423;
wire n_424;
wire n_897;
wire n_425;
wire n_426;
wire n_954;
wire n_427;
wire n_428;
wire n_1014;
wire n_429;
wire n_430;
wire n_1109;
wire n_431;
wire n_432;
wire n_1218;
wire n_433;
wire n_434;
wire n_1336;
wire n_435;
wire n_436;
wire n_1464;
wire n_437;
wire n_438;
wire n_1592;
wire n_439;
wire n_440;
wire n_1725;
wire n_441;
wire n_443;
wire n_442;
wire n_444;
wire n_1868;
wire n_2018;
wire n_445;
wire n_446;
wire n_2155;
wire n_448;
wire n_449;
wire n_450;
wire n_2644;
wire n_3509;
wire n_4205;
wire n_4563;
wire n_4655;
wire n_4762;
wire n_4873;
wire n_4951;
wire n_4956;
wire n_5118;
wire n_5159;
wire n_5238;
wire n_5368;
wire n_5426;
wire n_5465;
wire n_451;
wire n_5470;
wire n_5466;
wire n_5480;
wire n_452;
wire n_5483;
wire n_5481;
wire n_5495;
wire n_5477;
wire n_5496;
wire n_5478;
wire n_5745;
wire n_5743;
wire n_453;
wire n_5748;
wire n_458;
wire n_457;
wire n_455;
wire n_456;
wire n_473;
wire n_470;
wire n_471;
wire n_472;
wire n_469;
wire n_459;
wire n_485;
wire n_463;
wire n_464;
wire n_468;
wire n_466;
wire n_467;
wire n_499;
wire n_488;
wire n_489;
wire n_486;
wire n_482;
wire n_483;
wire n_478;
wire n_474;
wire n_475;
wire n_509;
wire n_477;
wire n_492;
wire n_480;
wire n_479;
wire n_481;
wire n_498;
wire n_487;
wire n_490;
wire n_503;
wire n_497;
wire n_496;
wire n_493;
wire n_525;
wire n_505;
wire n_501;
wire n_491;
wire n_506;
wire n_494;
wire n_495;
wire n_514;
wire n_515;
wire n_510;
wire n_500;
wire n_517;
wire n_502;
wire n_504;
wire n_531;
wire n_530;
wire n_526;
wire n_545;
wire n_523;
wire n_521;
wire n_507;
wire n_519;
wire n_512;
wire n_511;
wire n_513;
wire n_551;
wire n_516;
wire n_537;
wire n_518;
wire n_570;
wire n_520;
wire n_569;
wire n_567;
wire n_522;
wire n_544;
wire n_524;
wire n_528;
wire n_527;
wire n_554;
wire n_556;
wire n_552;
wire n_529;
wire n_5767;
wire n_5753;
wire n_532;
wire n_571;
wire n_549;
wire n_548;
wire n_542;
wire n_541;
wire n_538;
wire n_533;
wire n_534;
wire n_591;
wire n_536;
wire n_562;
wire n_539;
wire n_540;
wire n_579;
wire n_546;
wire n_566;
wire n_547;
wire n_563;
wire n_550;
wire n_553;
wire n_555;
wire n_557;
wire n_558;
wire n_575;
wire n_613;
wire n_580;
wire n_578;
wire n_576;
wire n_583;
wire n_585;
wire n_581;
wire n_559;
wire n_560;
wire n_625;
wire n_564;
wire n_565;
wire n_618;
wire n_617;
wire n_645;
wire n_619;
wire n_616;
wire n_568;
wire n_608;
wire n_572;
wire n_607;
wire n_573;
wire n_600;
wire n_574;
wire n_593;
wire n_611;
wire n_615;
wire n_609;
wire n_577;
wire n_612;
wire n_582;
wire n_584;
wire n_599;
wire n_586;
wire n_601;
wire n_606;
wire n_587;
wire n_604;
wire n_635;
wire n_598;
wire n_597;
wire n_594;
wire n_588;
wire n_589;
wire n_660;
wire n_592;
wire n_627;
wire n_595;
wire n_596;
wire n_657;
wire n_5750;
wire n_634;
wire n_630;
wire n_602;
wire n_638;
wire n_603;
wire n_629;
wire n_605;
wire n_610;
wire n_614;
wire n_644;
wire n_642;
wire n_640;
wire n_620;
wire n_646;
wire n_650;
wire n_652;
wire n_648;
wire n_656;
wire n_621;
wire n_655;
wire n_653;
wire n_622;
wire n_623;
wire n_701;
wire n_626;
wire n_675;
wire n_628;
wire n_661;
wire n_632;
wire n_631;
wire n_633;
wire n_685;
wire n_636;
wire n_684;
wire n_637;
wire n_672;
wire n_641;
wire n_643;
wire n_742;
wire n_721;
wire n_692;
wire n_690;
wire n_688;
wire n_647;
wire n_676;
wire n_649;
wire n_651;
wire n_691;
wire n_654;
wire n_668;
wire n_658;
wire n_667;
wire n_659;
wire n_680;
wire n_686;
wire n_687;
wire n_683;
wire n_666;
wire n_665;
wire n_662;
wire n_697;
wire n_695;
wire n_693;
wire n_663;
wire n_664;
wire n_737;
wire n_669;
wire n_670;
wire n_749;
wire n_673;
wire n_706;
wire n_674;
wire n_705;
wire n_677;
wire n_703;
wire n_678;
wire n_702;
wire n_679;
wire n_714;
wire n_733;
wire n_736;
wire n_731;
wire n_681;
wire n_682;
wire n_689;
wire n_720;
wire n_694;
wire n_696;
wire n_741;
wire n_710;
wire n_709;
wire n_707;
wire n_728;
wire n_730;
wire n_726;
wire n_719;
wire n_718;
wire n_715;
wire n_740;
wire n_744;
wire n_738;
wire n_698;
wire n_699;
wire n_794;
wire n_777;
wire n_704;
wire n_776;
wire n_774;
wire n_708;
wire n_787;
wire n_815;
wire n_788;
wire n_712;
wire n_711;
wire n_713;
wire n_751;
wire n_716;
wire n_717;
wire n_778;
wire n_722;
wire n_753;
wire n_723;
wire n_755;
wire n_724;
wire n_761;
wire n_725;
wire n_772;
wire n_727;
wire n_729;
wire n_767;
wire n_732;
wire n_734;
wire n_739;
wire n_743;
wire n_745;
wire n_771;
wire n_766;
wire n_762;
wire n_782;
wire n_784;
wire n_780;
wire n_758;
wire n_760;
wire n_756;
wire n_746;
wire n_747;
wire n_841;
wire n_750;
wire n_797;
wire n_752;
wire n_800;
wire n_754;
wire n_802;
wire n_757;
wire n_759;
wire n_835;
wire n_764;
wire n_763;
wire n_765;
wire n_825;
wire n_768;
wire n_824;
wire n_769;
wire n_795;
wire n_770;
wire n_811;
wire n_828;
wire n_830;
wire n_826;
wire n_773;
wire n_801;
wire n_775;
wire n_807;
wire n_779;
wire n_806;
wire n_781;
wire n_783;
wire n_785;
wire n_786;
wire n_5762;
wire n_789;
wire n_819;
wire n_823;
wire n_790;
wire n_821;
wire n_872;
wire n_805;
wire n_809;
wire n_808;
wire n_883;
wire n_836;
wire n_834;
wire n_832;
wire n_814;
wire n_816;
wire n_812;
wire n_791;
wire n_792;
wire n_898;
wire n_796;
wire n_845;
wire n_798;
wire n_853;
wire n_799;
wire n_844;
wire n_871;
wire n_867;
wire n_803;
wire n_804;
wire n_810;
wire n_842;
wire n_813;
wire n_817;
wire n_851;
wire n_5751;
wire n_818;
wire n_856;
wire n_881;
wire n_885;
wire n_879;
wire n_820;
wire n_865;
wire n_822;
wire n_827;
wire n_829;
wire n_833;
wire n_882;
wire n_888;
wire n_889;
wire n_886;
wire n_837;
wire n_843;
wire n_859;
wire n_861;
wire n_857;
wire n_876;
wire n_878;
wire n_874;
wire n_850;
wire n_849;
wire n_846;
wire n_838;
wire n_839;
wire n_955;
wire n_906;
wire n_907;
wire n_903;
wire n_847;
wire n_848;
wire n_949;
wire n_852;
wire n_901;
wire n_854;
wire n_913;
wire n_855;
wire n_899;
wire n_858;
wire n_860;
wire n_937;
wire n_862;
wire n_911;
wire n_863;
wire n_916;
wire n_864;
wire n_902;
wire n_866;
wire n_925;
wire n_869;
wire n_868;
wire n_870;
wire n_932;
wire n_873;
wire n_931;
wire n_875;
wire n_877;
wire n_908;
wire n_880;
wire n_884;
wire n_944;
wire n_887;
wire n_921;
wire n_919;
wire n_917;
wire n_890;
wire n_922;
wire n_891;
wire n_924;
wire n_892;
wire n_993;
wire n_929;
wire n_928;
wire n_936;
wire n_893;
wire n_935;
wire n_933;
wire n_941;
wire n_943;
wire n_939;
wire n_948;
wire n_894;
wire n_947;
wire n_945;
wire n_895;
wire n_896;
wire n_1015;
wire n_900;
wire n_966;
wire n_904;
wire n_905;
wire n_998;
wire n_909;
wire n_965;
wire n_910;
wire n_956;
wire n_912;
wire n_957;
wire n_914;
wire n_982;
wire n_915;
wire n_970;
wire n_918;
wire n_920;
wire n_1100;
wire n_923;
wire n_974;
wire n_1002;
wire n_1004;
wire n_1000;
wire n_992;
wire n_926;
wire n_990;
wire n_988;
wire n_930;
wire n_934;
wire n_964;
wire n_938;
wire n_963;
wire n_940;
wire n_942;
wire n_946;
wire n_980;
wire n_950;
wire n_971;
wire n_951;
wire n_986;
wire n_962;
wire n_961;
wire n_958;
wire n_1081;
wire n_999;
wire n_997;
wire n_995;
wire n_979;
wire n_978;
wire n_975;
wire n_1009;
wire n_1007;
wire n_1005;
wire n_952;
wire n_953;
wire n_1110;
wire n_959;
wire n_960;
wire n_1067;
wire n_967;
wire n_1026;
wire n_968;
wire n_1024;
wire n_969;
wire n_1016;
wire n_1088;
wire n_972;
wire n_1087;
wire n_1085;
wire n_973;
wire n_1025;
wire n_976;
wire n_977;
wire n_1089;
wire n_981;
wire n_1038;
wire n_983;
wire n_1041;
wire n_984;
wire n_1044;
wire n_985;
wire n_1017;
wire n_1066;
wire n_987;
wire n_1065;
wire n_1063;
wire n_989;
wire n_1023;
wire n_994;
wire n_1021;
wire n_996;
wire n_1080;
wire n_1001;
wire n_1003;
wire n_1054;
wire n_1006;
wire n_1008;
wire n_1096;
wire n_1032;
wire n_1031;
wire n_1027;
wire n_1010;
wire n_1060;
wire n_1011;
wire n_1181;
wire n_1019;
wire n_1018;
wire n_1079;
wire n_1083;
wire n_1075;
wire n_1051;
wire n_1050;
wire n_1047;
wire n_1095;
wire n_1094;
wire n_1090;
wire n_1012;
wire n_1013;
wire n_1222;
wire n_1020;
wire n_1028;
wire n_1204;
wire n_1279;
wire n_1208;
wire n_1035;
wire n_1033;
wire n_1036;
wire n_1116;
wire n_1037;
wire n_1119;
wire n_1193;
wire n_1042;
wire n_1191;
wire n_1189;
wire n_1043;
wire n_1134;
wire n_1048;
wire n_1049;
wire n_1194;
wire n_1055;
wire n_1142;
wire n_1057;
wire n_1117;
wire n_1058;
wire n_1120;
wire n_1059;
wire n_1144;
wire n_1180;
wire n_1061;
wire n_1177;
wire n_1172;
wire n_1062;
wire n_1155;
wire n_1064;
wire n_1152;
wire n_1071;
wire n_1151;
wire n_1076;
wire n_1082;
wire n_1187;
wire n_1086;
wire n_1129;
wire n_1091;
wire n_1093;
wire n_1201;
wire n_1104;
wire n_1162;
wire n_1105;
wire n_1143;
wire n_1150;
wire n_1149;
wire n_1145;
wire n_1298;
wire n_1188;
wire n_1185;
wire n_1183;
wire n_1125;
wire n_1124;
wire n_1121;
wire n_1198;
wire n_1200;
wire n_1196;
wire n_1108;
wire n_1115;
wire n_1111;
wire n_1112;
wire n_1346;
wire n_1118;
wire n_1236;
wire n_1122;
wire n_1123;
wire n_1319;
wire n_1138;
wire n_1234;
wire n_1139;
wire n_1226;
wire n_1140;
wire n_1228;
wire n_1405;
wire n_1292;
wire n_1290;
wire n_1288;
wire n_1146;
wire n_1148;
wire n_1291;
wire n_1153;
wire n_1231;
wire n_1156;
wire n_1284;
wire n_1157;
wire n_1265;
wire n_1158;
wire n_1248;
wire n_1309;
wire n_1318;
wire n_1304;
wire n_1167;
wire n_1285;
wire n_1176;
wire n_1259;
wire n_1182;
wire n_1255;
wire n_1184;
wire n_1297;
wire n_1190;
wire n_1247;
wire n_1195;
wire n_1246;
wire n_1197;
wire n_1199;
wire n_1202;
wire n_1203;
wire n_5758;
wire n_1209;
wire n_1233;
wire n_1263;
wire n_1264;
wire n_1254;
wire n_1295;
wire n_1300;
wire n_1293;
wire n_1243;
wire n_1242;
wire n_1237;
wire n_1329;
wire n_1332;
wire n_1324;
wire n_1278;
wire n_1277;
wire n_1269;
wire n_1212;
wire n_1213;
wire n_1465;
wire n_1223;
wire n_1340;
wire n_1225;
wire n_1337;
wire n_1227;
wire n_1353;
wire n_1229;
wire n_1350;
wire n_1230;
wire n_1342;
wire n_1377;
wire n_1381;
wire n_1371;
wire n_1235;
wire n_1356;
wire n_1240;
wire n_1241;
wire n_1413;
wire n_1249;
wire n_1250;
wire n_1273;
wire n_1274;
wire n_1430;
wire n_1280;
wire n_1347;
wire n_1281;
wire n_1367;
wire n_1360;
wire n_1363;
wire n_1357;
wire n_1286;
wire n_1393;
wire n_1287;
wire n_1354;
wire n_1289;
wire n_1404;
wire n_1294;
wire n_1299;
wire n_1305;
wire n_1314;
wire n_1328;
wire n_1331;
wire n_1361;
wire n_1455;
wire n_1450;
wire n_1434;
wire n_1333;
wire n_1392;
wire n_1397;
wire n_1399;
wire n_1395;
wire n_1403;
wire n_1409;
wire n_1401;
wire n_1557;
wire n_1414;
wire n_1412;
wire n_1410;
wire n_1418;
wire n_1421;
wire n_1416;
wire n_1424;
wire n_1426;
wire n_1422;
wire n_1334;
wire n_1335;
wire n_1577;
wire n_1339;
wire n_1470;
wire n_1341;
wire n_1481;
wire n_1343;
wire n_1471;
wire n_1348;
wire n_1496;
wire n_1349;
wire n_1466;
wire n_1352;
wire n_1483;
wire n_1355;
wire n_1533;
wire n_1358;
wire n_1362;
wire n_1564;
wire n_1372;
wire n_1373;
wire n_1551;
wire n_1382;
wire n_1493;
wire n_1387;
wire n_1491;
wire n_1388;
wire n_1472;
wire n_1391;
wire n_1501;
wire n_1512;
wire n_1517;
wire n_1502;
wire n_1486;
wire n_1488;
wire n_1484;
wire n_1396;
wire n_1398;
wire n_1542;
wire n_1402;
wire n_1406;
wire n_1411;
wire n_1556;
wire n_1417;
wire n_1419;
wire n_1521;
wire n_1423;
wire n_1425;
wire n_1440;
wire n_1435;
wire n_1478;
wire n_1475;
wire n_1473;
wire n_1445;
wire n_5757;
wire n_1459;
wire n_1535;
wire n_1541;
wire n_1460;
wire n_1539;
wire n_1537;
wire n_1546;
wire n_1550;
wire n_1544;
wire n_1554;
wire n_1559;
wire n_1552;
wire n_1631;
wire n_1565;
wire n_1563;
wire n_1560;
wire n_1568;
wire n_1570;
wire n_1566;
wire n_1462;
wire n_1463;
wire n_1721;
wire n_1467;
wire n_1598;
wire n_1474;
wire n_1477;
wire n_1714;
wire n_1479;
wire n_1597;
wire n_1480;
wire n_1582;
wire n_1485;
wire n_1487;
wire n_1490;
wire n_1607;
wire n_1492;
wire n_1611;
wire n_1497;
wire n_1649;
wire n_1506;
wire n_1507;
wire n_1703;
wire n_1522;
wire n_1622;
wire n_1527;
wire n_1583;
wire n_1531;
wire n_1634;
wire n_1532;
wire n_1625;
wire n_1629;
wire n_1633;
wire n_1626;
wire n_1615;
wire n_1617;
wire n_1612;
wire n_1536;
wire n_1638;
wire n_1538;
wire n_1658;
wire n_1543;
wire n_1657;
wire n_1545;
wire n_1549;
wire n_1553;
wire n_1558;
wire n_1692;
wire n_1562;
wire n_1630;
wire n_1567;
wire n_1569;
wire n_1707;
wire n_1571;
wire n_1623;
wire n_1572;
wire n_1646;
wire n_1653;
wire n_1573;
wire n_1651;
wire n_1811;
wire n_1668;
wire n_1672;
wire n_1662;
wire n_1683;
wire n_1687;
wire n_1677;
wire n_1700;
wire n_1702;
wire n_1696;
wire n_1706;
wire n_1709;
wire n_1704;
wire n_1853;
wire n_1716;
wire n_1710;
wire n_1586;
wire n_1791;
wire n_1587;
wire n_1591;
wire n_1872;
wire n_1601;
wire n_1756;
wire n_1602;
wire n_1726;
wire n_1613;
wire n_1616;
wire n_1785;
wire n_1618;
wire n_1729;
wire n_1619;
wire n_1734;
wire n_1919;
wire n_1839;
wire n_1834;
wire n_1832;
wire n_1624;
wire n_1727;
wire n_1628;
wire n_1632;
wire n_1636;
wire n_1803;
wire n_1637;
wire n_1730;
wire n_1639;
wire n_1640;
wire n_1798;
wire n_1793;
wire n_1796;
wire n_1797;
wire n_1792;
wire n_1643;
wire n_1786;
wire n_1644;
wire n_1735;
wire n_1645;
wire n_1766;
wire n_1822;
wire n_1824;
wire n_1820;
wire n_1810;
wire n_1650;
wire n_1807;
wire n_1805;
wire n_1652;
wire n_1667;
wire n_1671;
wire n_1682;
wire n_1686;
wire n_1697;
wire n_1701;
wire n_1705;
wire n_1708;
wire n_1838;
wire n_1711;
wire n_1715;
wire n_1717;
wire n_1731;
wire n_1718;
wire n_1801;
wire n_1817;
wire n_1819;
wire n_1813;
wire n_1781;
wire n_1776;
wire n_1767;
wire n_1827;
wire n_1831;
wire n_1825;
wire n_1741;
wire n_1746;
wire n_1745;
wire n_2003;
wire n_1847;
wire n_1843;
wire n_1722;
wire n_1882;
wire n_1723;
wire n_1724;
wire n_2019;
wire n_1728;
wire n_1906;
wire n_1732;
wire n_2056;
wire n_1997;
wire n_1996;
wire n_1992;
wire n_1736;
wire n_1737;
wire n_1747;
wire n_1893;
wire n_1750;
wire n_1895;
wire n_1751;
wire n_1883;
wire n_1757;
wire n_1910;
wire n_1761;
wire n_1902;
wire n_1771;
wire n_1775;
wire n_1789;
wire n_1903;
wire n_1790;
wire n_1908;
wire n_2009;
wire n_2010;
wire n_2006;
wire n_1799;
wire n_1921;
wire n_1800;
wire n_1885;
wire n_1802;
wire n_2070;
wire n_1985;
wire n_1984;
wire n_1975;
wire n_1804;
wire n_1950;
wire n_1806;
wire n_1890;
wire n_1812;
wire n_1889;
wire n_1814;
wire n_1818;
wire n_1821;
wire n_1823;
wire n_1929;
wire n_1826;
wire n_1828;
wire n_1833;
wire n_1918;
wire n_1844;
wire n_2002;
wire n_1848;
wire n_1858;
wire n_1945;
wire n_1862;
wire n_1907;
wire n_1863;
wire n_2108;
wire n_1887;
wire n_1886;
wire n_1965;
wire n_1974;
wire n_1960;
wire n_1928;
wire n_1927;
wire n_1922;
wire n_1989;
wire n_1991;
wire n_1986;
wire n_1917;
wire n_1916;
wire n_1911;
wire n_2001;
wire n_2005;
wire n_1998;
wire n_1864;
wire n_1878;
wire n_1873;
wire n_1898;
wire n_1888;
wire n_1894;
wire n_2028;
wire n_1896;
wire n_1897;
wire n_2210;
wire n_1900;
wire n_2023;
wire n_1901;
wire n_2025;
wire n_1904;
wire n_2035;
wire n_2118;
wire n_2122;
wire n_2116;
wire n_1909;
wire n_2042;
wire n_1914;
wire n_1915;
wire n_2136;
wire n_1923;
wire n_1924;
wire n_2123;
wire n_1930;
wire n_2032;
wire n_1931;
wire n_2036;
wire n_1935;
wire n_2029;
wire n_1939;
wire n_2086;
wire n_1940;
wire n_2057;
wire n_2132;
wire n_2135;
wire n_2130;
wire n_2106;
wire n_1954;
wire n_2105;
wire n_2103;
wire n_1955;
wire n_2080;
wire n_1964;
wire n_1970;
wire n_2114;
wire n_1980;
wire n_1988;
wire n_1990;
wire n_1995;
wire n_1999;
wire n_2004;
wire n_2007;
wire n_2011;
wire n_2096;
wire n_2012;
wire n_2101;
wire n_2013;
wire n_2102;
wire n_2233;
wire n_2115;
wire n_2112;
wire n_2110;
wire n_2258;
wire n_2066;
wire n_2060;
wire n_2126;
wire n_2129;
wire n_2124;
wire n_2284;
wire n_2055;
wire n_2045;
wire n_2139;
wire n_2143;
wire n_2137;
wire n_2094;
wire n_2095;
wire n_2090;
wire n_2016;
wire n_2017;
wire n_2334;
wire n_2020;
wire n_2161;
wire n_2022;
wire n_2159;
wire n_2024;
wire n_2180;
wire n_2026;
wire n_2204;
wire n_2027;
wire n_2170;
wire n_2030;
wire n_2235;
wire n_2031;
wire n_2174;
wire n_2460;
wire n_2195;
wire n_2190;
wire n_2185;
wire n_2041;
wire n_2184;
wire n_2046;
wire n_2051;
wire n_2061;
wire n_2062;
wire n_2071;
wire n_2213;
wire n_2076;
wire n_2208;
wire n_2081;
wire n_2240;
wire n_2091;
wire n_2093;
wire n_2309;
wire n_2097;
wire n_2215;
wire n_2098;
wire n_2224;
wire n_2219;
wire n_2222;
wire n_2216;
wire n_2230;
wire n_2231;
wire n_2225;
wire n_2104;
wire n_2247;
wire n_2109;
wire n_2246;
wire n_2111;
wire n_2232;
wire n_2117;
wire n_2119;
wire n_2125;
wire n_2127;
wire n_2223;
wire n_2131;
wire n_2133;
wire n_2138;
wire n_2140;
wire n_2325;
wire n_2324;
wire n_2313;
wire n_2144;
wire n_2239;
wire n_2145;
wire n_2214;
wire n_2245;
wire n_2252;
wire n_2251;
wire n_2446;
wire n_2256;
wire n_2253;
wire n_2264;
wire n_2268;
wire n_2259;
wire n_2146;
wire n_2456;
wire n_2279;
wire n_2269;
wire n_2289;
wire n_2299;
wire n_2285;
wire n_2466;
wire n_2304;
wire n_2300;
wire n_2150;
wire n_2154;
wire n_2474;
wire n_2160;
wire n_2338;
wire n_2165;
wire n_2335;
wire n_2171;
wire n_2345;
wire n_2175;
wire n_2362;
wire n_2186;
wire n_2194;
wire n_2200;
wire n_2343;
wire n_2205;
wire n_2358;
wire n_2209;
wire n_2375;
wire n_2211;
wire n_2363;
wire n_2212;
wire n_2355;
wire n_2391;
wire n_2382;
wire n_2376;
wire n_2217;
wire n_2218;
wire n_2226;
wire n_2229;
wire n_2234;
wire n_2336;
wire n_2236;
wire n_2412;
wire n_2237;
wire n_2346;
wire n_2238;
wire n_2369;
wire n_2349;
wire n_2524;
wire n_2350;
wire n_2372;
wire n_2548;
wire n_2371;
wire n_2243;
wire n_2397;
wire n_2244;
wire n_2250;
wire n_2254;
wire n_2257;
wire n_2260;
wire n_2265;
wire n_2373;
wire n_2274;
wire n_2288;
wire n_2294;
wire n_2351;
wire n_2303;
wire n_2305;
wire n_2319;
wire n_2314;
wire n_2367;
wire n_2487;
wire n_2365;
wire n_2323;
wire n_5756;
wire n_2326;
wire n_2359;
wire n_2327;
wire n_2417;
wire n_2427;
wire n_2585;
wire n_2432;
wire n_2437;
wire n_2328;
wire n_2590;
wire n_2442;
wire n_2450;
wire n_2603;
wire n_2452;
wire n_2454;
wire n_2329;
wire n_2607;
wire n_2455;
wire n_2458;
wire n_2330;
wire n_2618;
wire n_2459;
wire n_2481;
wire n_2625;
wire n_2464;
wire n_2331;
wire n_2472;
wire n_2337;
wire n_2527;
wire n_2341;
wire n_2475;
wire n_2342;
wire n_2477;
wire n_2344;
wire n_2497;
wire n_2523;
wire n_2347;
wire n_2348;
wire n_2352;
wire n_2489;
wire n_2356;
wire n_2492;
wire n_2357;
wire n_2478;
wire n_2598;
wire n_2599;
wire n_2595;
wire n_2364;
wire n_2366;
wire n_5755;
wire n_2368;
wire n_2500;
wire n_2547;
wire n_2370;
wire n_2594;
wire n_2378;
wire n_2377;
wire n_2387;
wire n_2392;
wire n_2506;
wire n_2402;
wire n_2493;
wire n_2406;
wire n_2479;
wire n_2407;
wire n_2509;
wire n_2408;
wire n_2498;
wire n_2617;
wire n_2616;
wire n_2612;
wire n_2583;
wire n_2582;
wire n_2577;
wire n_2422;
wire n_2501;
wire n_2584;
wire n_2426;
wire n_2428;
wire n_2436;
wire n_2528;
wire n_2602;
wire n_2447;
wire n_2451;
wire n_2610;
wire n_2453;
wire n_2513;
wire n_2457;
wire n_2619;
wire n_2624;
wire n_2461;
wire n_2480;
wire n_2465;
wire n_2638;
wire n_2631;
wire n_2467;
wire n_2567;
wire n_2468;
wire n_2568;
wire n_2589;
wire n_2592;
wire n_2586;
wire n_2543;
wire n_2539;
wire n_2606;
wire n_2611;
wire n_2609;
wire n_2522;
wire n_2518;
wire n_2623;
wire n_2627;
wire n_2471;
wire n_2819;
wire n_2485;
wire n_2473;
wire n_2649;
wire n_2476;
wire n_2699;
wire n_2482;
wire n_2486;
wire n_2488;
wire n_2658;
wire n_2765;
wire n_2494;
wire n_2763;
wire n_2761;
wire n_2495;
wire n_2650;
wire n_2496;
wire n_2669;
wire n_2749;
wire n_2499;
wire n_2502;
wire n_2674;
wire n_2503;
wire n_2675;
wire n_2507;
wire n_2726;
wire n_2508;
wire n_2704;
wire n_2514;
wire n_2517;
wire n_2779;
wire n_2533;
wire n_2538;
wire n_2766;
wire n_2553;
wire n_2673;
wire n_2557;
wire n_2714;
wire n_2558;
wire n_2733;
wire n_2559;
wire n_2719;
wire n_2563;
wire n_2679;
wire n_2872;
wire n_2780;
wire n_2778;
wire n_2774;
wire n_2752;
wire n_2748;
wire n_2745;
wire n_2573;
wire n_2738;
wire n_2578;
wire n_2581;
wire n_2760;
wire n_2588;
wire n_2591;
wire n_2596;
wire n_2597;
wire n_2773;
wire n_2604;
wire n_2605;
wire n_2613;
wire n_2615;
wire n_2800;
wire n_2620;
wire n_2626;
wire n_2628;
wire n_2632;
wire n_2630;
wire n_2637;
wire n_2633;
wire n_2813;
wire n_2636;
wire n_2814;
wire n_2804;
wire n_5754;
wire n_2639;
wire n_2830;
wire n_2833;
wire n_2824;
wire n_2640;
wire n_2742;
wire n_2643;
wire n_2744;
wire n_2755;
wire n_2759;
wire n_2753;
wire n_2695;
wire n_2694;
wire n_2684;
wire n_2770;
wire n_2772;
wire n_2768;
wire n_2732;
wire n_2731;
wire n_2727;
wire n_2794;
wire n_2799;
wire n_2784;
wire n_2725;
wire n_2724;
wire n_2720;
wire n_2654;
wire n_2857;
wire n_2655;
wire n_2839;
wire n_2659;
wire n_2860;
wire n_2660;
wire n_2843;
wire n_2664;
wire n_2853;
wire n_2870;
wire n_2874;
wire n_2867;
wire n_2689;
wire n_2693;
wire n_2962;
wire n_2703;
wire n_2861;
wire n_2709;
wire n_2858;
wire n_2713;
wire n_2865;
wire n_2717;
wire n_2866;
wire n_2718;
wire n_2880;
wire n_2721;
wire n_2723;
wire n_3013;
wire n_2728;
wire n_2729;
wire n_2997;
wire n_2734;
wire n_2923;
wire n_2735;
wire n_2878;
wire n_2917;
wire n_2916;
wire n_2914;
wire n_2739;
wire n_2881;
wire n_2740;
wire n_2892;
wire n_2741;
wire n_2901;
wire n_2896;
wire n_2897;
wire n_2893;
wire n_3106;
wire n_2908;
wire n_2906;
wire n_2902;
wire n_2747;
wire n_2746;
wire n_2750;
wire n_2754;
wire n_2756;
wire n_2762;
wire n_2900;
wire n_2767;
wire n_2899;
wire n_2769;
wire n_2771;
wire n_2775;
wire n_2871;
wire n_2789;
wire n_2798;
wire n_2809;
wire n_2889;
wire n_2825;
wire n_2888;
wire n_2887;
wire n_2882;
wire n_2829;
wire n_2834;
wire n_2922;
wire n_2835;
wire n_2879;
wire n_2936;
wire n_2942;
wire n_2932;
wire n_2951;
wire n_2957;
wire n_2947;
wire n_2972;
wire n_2978;
wire n_2963;
wire n_2992;
wire n_2987;
wire n_2981;
wire n_3003;
wire n_3005;
wire n_3001;
wire n_3008;
wire n_3012;
wire n_3006;
wire n_2844;
wire n_3024;
wire n_2849;
wire n_3020;
wire n_2854;
wire n_3036;
wire n_2855;
wire n_3021;
wire n_2859;
wire n_3063;
wire n_2864;
wire n_3050;
wire n_2868;
wire n_2873;
wire n_3163;
wire n_2875;
wire n_3041;
wire n_2876;
wire n_3025;
wire n_3120;
wire n_3125;
wire n_3114;
wire n_2885;
wire n_2886;
wire n_3258;
wire n_2891;
wire n_3037;
wire n_2894;
wire n_2895;
wire n_3141;
wire n_2903;
wire n_3105;
wire n_2907;
wire n_2909;
wire n_3047;
wire n_2910;
wire n_3042;
wire n_2912;
wire n_3026;
wire n_2913;
wire n_3054;
wire n_2915;
wire n_2921;
wire n_2920;
wire n_3168;
wire n_3171;
wire n_3166;
wire n_3174;
wire n_3176;
wire n_3172;
wire n_3154;
wire n_3158;
wire n_3145;
wire n_2926;
wire n_3051;
wire n_2927;
wire n_3071;
wire n_2933;
wire n_2937;
wire n_3069;
wire n_2948;
wire n_2952;
wire n_2967;
wire n_2977;
wire n_3062;
wire n_2982;
wire n_2991;
wire n_3002;
wire n_3004;
wire n_3034;
wire n_3007;
wire n_3009;
wire n_3014;
wire n_3085;
wire n_3015;
wire n_3090;
wire n_3100;
wire n_3111;
wire n_3095;
wire n_3068;
wire n_3067;
wire n_3064;
wire n_3140;
wire n_3016;
wire n_3135;
wire n_3130;
wire n_3061;
wire n_3058;
wire n_3055;
wire n_3162;
wire n_3019;
wire n_3161;
wire n_3159;
wire n_3033;
wire n_3030;
wire n_3027;
wire n_3022;
wire n_3188;
wire n_3023;
wire n_3181;
wire n_3028;
wire n_3029;
wire n_3330;
wire n_3035;
wire n_3182;
wire n_3040;
wire n_3210;
wire n_3043;
wire n_3246;
wire n_3044;
wire n_3183;
wire n_3045;
wire n_3202;
wire n_3046;
wire n_3189;
wire n_3048;
wire n_3223;
wire n_3049;
wire n_3207;
wire n_3364;
wire n_3238;
wire n_3236;
wire n_3227;
wire n_3056;
wire n_3057;
wire n_3315;
wire n_3065;
wire n_3066;
wire n_3293;
wire n_3070;
wire n_3203;
wire n_3075;
wire n_3403;
wire n_3252;
wire n_3247;
wire n_3079;
wire n_3214;
wire n_3080;
wire n_3190;
wire n_3217;
wire n_3220;
wire n_3215;
wire n_3200;
wire n_3195;
wire n_3192;
wire n_3091;
wire n_3271;
wire n_3099;
wire n_3110;
wire n_3237;
wire n_3115;
wire n_3124;
wire n_3302;
wire n_3134;
wire n_3197;
wire n_3144;
wire n_3196;
wire n_3150;
wire n_3155;
wire n_3322;
wire n_3160;
wire n_3222;
wire n_3165;
wire n_3221;
wire n_3167;
wire n_3169;
wire n_3173;
wire n_3175;
wire n_3179;
wire n_3267;
wire n_3180;
wire n_3211;
wire n_3282;
wire n_3292;
wire n_3277;
wire n_3301;
wire n_3311;
wire n_3297;
wire n_3466;
wire n_3316;
wire n_3314;
wire n_3312;
wire n_3319;
wire n_3324;
wire n_3317;
wire n_3488;
wire n_3331;
wire n_3329;
wire n_3325;
wire n_3336;
wire n_3334;
wire n_3332;
wire n_3184;
wire n_3352;
wire n_3186;
wire n_3339;
wire n_3187;
wire n_3340;
wire n_3193;
wire n_3194;
wire n_3201;
wire n_3347;
wire n_3204;
wire n_3381;
wire n_3205;
wire n_3343;
wire n_3208;
wire n_3373;
wire n_3209;
wire n_3354;
wire n_3545;
wire n_3452;
wire n_3443;
wire n_3441;
wire n_3213;
wire n_3365;
wire n_3216;
wire n_3218;
wire n_3232;
wire n_3361;
wire n_3242;
wire n_3368;
wire n_3496;
wire n_3495;
wire n_3491;
wire n_3257;
wire n_3262;
wire n_3375;
wire n_3263;
wire n_3355;
wire n_3526;
wire n_3481;
wire n_3479;
wire n_3476;
wire n_3272;
wire n_3417;
wire n_3276;
wire n_3366;
wire n_3281;
wire n_3287;
wire n_3298;
wire n_3307;
wire n_3447;
wire n_3313;
wire n_3462;
wire n_3318;
wire n_3323;
wire n_3480;
wire n_3326;
wire n_3485;
wire n_3333;
wire n_3335;
wire n_3497;
wire n_3337;
wire n_3412;
wire n_3411;
wire n_3407;
wire n_3338;
wire n_3371;
wire n_3360;
wire n_3359;
wire n_3356;
wire n_3432;
wire n_3437;
wire n_3427;
wire n_3385;
wire n_3387;
wire n_3382;
wire n_3458;
wire n_3472;
wire n_3453;
wire n_3380;
wire n_3379;
wire n_3376;
wire n_3484;
wire n_3490;
wire n_3482;
wire n_3344;
wire n_3517;
wire n_3345;
wire n_3501;
wire n_3346;
wire n_3502;
wire n_3350;
wire n_3503;
wire n_3351;
wire n_3512;
wire n_3353;
wire n_3527;
wire n_3357;
wire n_3358;
wire n_3597;
wire n_3367;
wire n_3505;
wire n_3644;
wire n_3372;
wire n_3643;
wire n_3638;
wire n_3374;
wire n_3518;
wire n_3377;
wire n_3378;
wire n_3655;
wire n_3384;
wire n_3386;
wire n_3637;
wire n_3388;
wire n_3504;
wire n_3392;
wire n_3533;
wire n_3396;
wire n_3546;
wire n_3397;
wire n_3551;
wire n_3402;
wire n_3537;
wire n_3406;
wire n_3679;
wire n_3662;
wire n_3659;
wire n_3657;
wire n_3413;
wire n_3554;
wire n_3558;
wire n_3552;
wire n_3608;
wire n_3618;
wire n_3598;
wire n_3422;
wire n_3573;
wire n_3431;
wire n_3433;
wire n_3442;
wire n_3544;
wire n_3457;
wire n_3467;
wire n_3647;
wire n_3478;
wire n_3525;
wire n_3483;
wire n_3489;
wire n_3492;
wire n_3493;
wire n_3498;
wire n_3568;
wire n_3587;
wire n_3593;
wire n_3583;
wire n_3543;
wire n_3541;
wire n_3538;
wire n_3627;
wire n_3633;
wire n_3619;
wire n_3524;
wire n_3523;
wire n_3519;
wire n_3654;
wire n_3499;
wire n_3652;
wire n_3650;
wire n_3902;
wire n_3766;
wire n_3764;
wire n_3759;
wire n_3506;
wire n_3511;
wire n_3510;
wire n_3514;
wire n_3513;
wire n_3531;
wire n_3516;
wire n_3667;
wire n_3520;
wire n_3522;
wire n_3765;
wire n_3530;
wire n_3665;
wire n_3532;
wire n_3671;
wire n_3534;
wire n_3672;
wire n_3535;
wire n_3684;
wire n_3539;
wire n_3540;
wire n_3740;
wire n_3547;
wire n_3711;
wire n_3548;
wire n_3687;
wire n_3553;
wire n_3557;
wire n_3806;
wire n_3559;
wire n_3691;
wire n_3563;
wire n_3700;
wire n_3731;
wire n_3739;
wire n_3729;
wire n_3578;
wire n_3715;
wire n_3584;
wire n_3588;
wire n_3603;
wire n_3613;
wire n_3706;
wire n_3623;
wire n_3628;
wire n_3639;
wire n_3699;
wire n_3648;
wire n_3698;
wire n_3651;
wire n_3784;
wire n_3656;
wire n_3781;
wire n_3658;
wire n_3680;
wire n_3663;
wire n_3796;
wire n_3800;
wire n_3794;
wire n_3664;
wire n_3841;
wire n_3840;
wire n_3837;
wire n_3720;
wire n_3725;
wire n_3718;
wire n_3705;
wire n_3708;
wire n_3701;
wire n_3750;
wire n_3756;
wire n_3744;
wire n_3697;
wire n_3696;
wire n_3692;
wire n_3780;
wire n_3790;
wire n_3770;
wire n_3678;
wire n_3677;
wire n_3673;
wire n_3666;
wire n_3817;
wire n_3669;
wire n_3819;
wire n_3670;
wire n_3818;
wire n_3675;
wire n_3676;
wire n_3683;
wire n_3831;
wire n_3685;
wire n_3847;
wire n_3686;
wire n_3833;
wire n_3688;
wire n_3821;
wire n_3690;
wire n_3820;
wire n_3693;
wire n_3694;
wire n_3704;
wire n_3707;
wire n_3709;
wire n_3844;
wire n_3712;
wire n_3868;
wire n_3713;
wire n_3836;
wire n_3714;
wire n_3851;
wire n_3854;
wire n_3858;
wire n_3852;
wire n_3719;
wire n_3721;
wire n_3730;
wire n_3735;
wire n_3745;
wire n_3755;
wire n_3760;
wire n_3897;
wire n_3775;
wire n_3785;
wire n_3917;
wire n_3795;
wire n_3805;
wire n_3826;
wire n_3825;
wire n_3822;
wire n_3810;
wire n_3866;
wire n_3865;
wire n_3864;
wire n_3862;
wire n_3815;
wire n_3850;
wire n_3874;
wire n_3878;
wire n_3872;
wire n_3881;
wire n_3883;
wire n_3879;
wire n_3886;
wire n_3888;
wire n_3884;
wire n_3896;
wire n_3911;
wire n_3892;
wire n_3995;
wire n_3922;
wire n_3916;
wire n_3912;
wire n_3823;
wire n_3824;
wire n_4146;
wire n_3829;
wire n_3933;
wire n_3830;
wire n_3936;
wire n_3832;
wire n_3937;
wire n_3838;
wire n_3839;
wire n_4032;
wire n_3842;
wire n_3952;
wire n_3843;
wire n_3957;
wire n_3845;
wire n_3958;
wire n_3846;
wire n_3982;
wire n_3968;
wire n_3973;
wire n_3962;
wire n_3853;
wire n_3857;
wire n_4018;
wire n_3859;
wire n_3976;
wire n_3860;
wire n_3988;
wire n_3861;
wire n_3996;
wire n_3863;
wire n_4045;
wire n_4041;
wire n_4039;
wire n_3867;
wire n_3993;
wire n_3992;
wire n_3989;
wire n_4003;
wire n_4000;
wire n_3997;
wire n_3871;
wire n_3984;
wire n_3873;
wire n_3875;
wire n_3880;
wire n_3882;
wire n_3885;
wire n_3887;
wire n_4004;
wire n_3893;
wire n_3907;
wire n_3913;
wire n_3994;
wire n_3927;
wire n_4011;
wire n_3928;
wire n_4012;
wire n_4015;
wire n_4017;
wire n_4013;
wire n_4021;
wire n_4025;
wire n_4019;
wire n_4031;
wire n_3932;
wire n_4028;
wire n_4026;
wire n_4036;
wire n_4038;
wire n_4034;
wire n_3942;
wire n_4069;
wire n_3943;
wire n_4048;
wire n_3947;
wire n_4049;
wire n_3953;
wire n_4052;
wire n_3956;
wire n_4064;
wire n_3967;
wire n_3972;
wire n_3977;
wire n_4110;
wire n_3987;
wire n_4152;
wire n_3990;
wire n_3991;
wire n_4186;
wire n_3998;
wire n_3999;
wire n_4173;
wire n_4005;
wire n_4053;
wire n_4006;
wire n_4075;
wire n_4007;
wire n_4134;
wire n_4010;
wire n_4080;
wire n_4099;
wire n_4104;
wire n_4084;
wire n_4119;
wire n_4129;
wire n_4114;
wire n_4014;
wire n_4016;
wire n_4020;
wire n_4024;
wire n_4027;
wire n_4109;
wire n_4033;
wire n_4105;
wire n_4035;
wire n_4037;
wire n_4179;
wire n_4040;
wire n_4042;
wire n_4046;
wire n_4054;
wire n_4158;
wire n_4160;
wire n_4154;
wire n_4163;
wire n_4166;
wire n_4161;
wire n_4169;
wire n_4172;
wire n_4167;
wire n_4203;
wire n_4180;
wire n_4176;
wire n_4174;
wire n_4184;
wire n_4047;
wire n_4183;
wire n_4181;
wire n_4304;
wire n_4306;
wire n_4301;
wire n_4055;
wire n_4190;
wire n_4059;
wire n_4192;
wire n_4065;
wire n_4193;
wire n_4068;
wire n_4207;
wire n_4074;
wire n_4268;
wire n_4078;
wire n_4194;
wire n_4079;
wire n_4238;
wire n_4089;
wire n_4094;
wire n_4324;
wire n_4115;
wire n_4124;
wire n_4312;
wire n_4130;
wire n_4208;
wire n_4138;
wire n_4149;
wire n_4148;
wire n_4139;
wire n_4144;
wire n_4283;
wire n_4150;
wire n_4330;
wire n_4333;
wire n_4327;
wire n_4151;
wire n_4247;
wire n_4318;
wire n_4320;
wire n_4315;
wire n_4153;
wire n_4269;
wire n_4155;
wire n_4159;
wire n_4162;
wire n_4165;
wire n_4264;
wire n_4168;
wire n_4171;
wire n_4175;
wire n_4202;
wire n_4182;
wire n_4335;
wire n_4187;
wire n_4334;
wire n_4188;
wire n_4292;
wire n_4289;
wire n_4288;
wire n_4189;
wire n_4298;
wire n_4309;
wire n_4314;
wire n_4307;
wire n_4263;
wire n_4262;
wire n_4248;
wire n_4438;
wire n_4326;
wire n_4323;
wire n_4321;
wire n_4201;
wire n_4200;
wire n_4195;
wire n_4196;
wire n_4197;
wire n_4452;
wire n_4204;
wire n_4213;
wire n_4209;
wire n_4228;
wire n_4212;
wire n_4223;
wire n_4214;
wire n_4343;
wire n_4218;
wire n_4337;
wire n_4233;
wire n_4341;
wire n_4504;
wire n_4340;
wire n_4239;
wire n_4344;
wire n_4243;
wire n_4350;
wire n_4253;
wire n_4258;
wire n_4417;
wire n_4273;
wire n_4383;
wire n_4278;
wire n_4351;
wire n_4282;
wire n_4360;
wire n_4284;
wire n_4479;
wire n_4450;
wire n_4443;
wire n_4293;
wire n_4356;
wire n_4359;
wire n_4354;
wire n_4413;
wire n_4300;
wire n_4408;
wire n_4403;
wire n_4303;
wire n_4305;
wire n_4308;
wire n_4313;
wire n_4316;
wire n_4319;
wire n_4372;
wire n_4322;
wire n_4434;
wire n_4328;
wire n_4329;
wire n_4543;
wire n_4336;
wire n_4345;
wire n_4339;
wire n_4393;
wire n_4398;
wire n_4388;
wire n_4368;
wire n_4364;
wire n_4361;
wire n_4433;
wire n_4442;
wire n_4423;
wire n_4342;
wire n_4456;
wire n_4512;
wire n_4514;
wire n_4510;
wire n_4347;
wire n_4457;
wire n_4348;
wire n_4466;
wire n_4349;
wire n_4458;
wire n_4355;
wire n_4357;
wire n_4362;
wire n_4363;
wire n_4517;
wire n_4373;
wire n_4459;
wire n_4378;
wire n_4470;
wire n_4379;
wire n_4472;
wire n_4382;
wire n_4483;
wire n_4499;
wire n_4501;
wire n_4497;
wire n_4384;
wire n_4462;
wire n_4389;
wire n_4397;
wire n_4404;
wire n_4488;
wire n_4418;
wire n_4487;
wire n_4428;
wire n_4439;
wire n_4448;
wire n_4480;
wire n_4453;
wire n_4454;
wire n_4614;
wire n_4537;
wire n_4534;
wire n_4455;
wire n_4496;
wire n_4507;
wire n_4509;
wire n_4505;
wire n_4486;
wire n_4491;
wire n_4490;
wire n_4528;
wire n_4533;
wire n_4518;
wire n_4478;
wire n_4477;
wire n_4473;
wire n_4463;
wire n_4622;
wire n_4464;
wire n_4552;
wire n_4465;
wire n_4553;
wire n_4467;
wire n_4558;
wire n_4469;
wire n_4568;
wire n_4471;
wire n_4607;
wire n_4475;
wire n_4476;
wire n_4611;
wire n_4484;
wire n_4485;
wire n_4492;
wire n_4600;
wire n_4493;
wire n_4602;
wire n_4494;
wire n_4573;
wire n_4588;
wire n_4587;
wire n_4578;
wire n_4498;
wire n_4500;
wire n_4506;
wire n_4508;
wire n_4635;
wire n_4511;
wire n_4513;
wire n_4523;
wire n_4529;
wire n_4650;
wire n_4758;
wire n_4612;
wire n_4610;
wire n_4608;
wire n_4538;
wire n_4616;
wire n_4548;
wire n_4617;
wire n_4625;
wire n_4629;
wire n_4623;
wire n_4632;
wire n_4634;
wire n_4630;
wire n_4638;
wire n_4642;
wire n_4636;
wire n_4645;
wire n_4649;
wire n_4643;
wire n_4559;
wire n_4694;
wire n_4562;
wire n_4598;
wire n_4583;
wire n_4584;
wire n_4743;
wire n_4593;
wire n_4595;
wire n_4765;
wire n_4599;
wire n_4660;
wire n_4601;
wire n_4705;
wire n_4603;
wire n_4700;
wire n_4604;
wire n_4699;
wire n_4609;
wire n_4755;
wire n_4613;
wire n_4665;
wire n_4615;
wire n_4621;
wire n_4618;
wire n_4675;
wire n_4680;
wire n_4666;
wire n_4754;
wire n_4760;
wire n_4752;
wire n_4715;
wire n_4721;
wire n_4709;
wire n_4624;
wire n_4628;
wire n_4631;
wire n_4633;
wire n_4637;
wire n_4639;
wire n_4644;
wire n_4646;
wire n_4651;
wire n_4730;
wire n_4737;
wire n_4739;
wire n_4735;
wire n_4838;
wire n_4744;
wire n_4742;
wire n_4740;
wire n_4747;
wire n_4751;
wire n_4745;
wire n_4654;
wire n_4690;
wire n_4670;
wire n_4679;
wire n_4853;
wire n_4681;
wire n_4685;
wire n_4874;
wire n_4695;
wire n_4779;
wire n_4701;
wire n_4807;
wire n_4710;
wire n_4720;
wire n_4818;
wire n_4724;
wire n_4775;
wire n_4725;
wire n_4766;
wire n_4833;
wire n_4842;
wire n_4828;
wire n_4732;
wire n_4789;
wire n_4736;
wire n_4738;
wire n_4772;
wire n_4741;
wire n_4834;
wire n_4746;
wire n_4748;
wire n_4785;
wire n_4753;
wire n_4759;
wire n_4870;
wire n_4865;
wire n_4868;
wire n_4858;
wire n_4769;
wire n_4774;
wire n_4767;
wire n_4817;
wire n_4823;
wire n_4808;
wire n_4784;
wire n_4783;
wire n_4780;
wire n_4849;
wire n_4857;
wire n_4843;
wire n_4761;
wire n_4764;
wire n_4763;
wire n_4787;
wire n_4768;
wire n_4773;
wire n_4776;
wire n_4886;
wire n_4781;
wire n_4782;
wire n_4894;
wire n_4786;
wire n_4793;
wire n_4788;
wire n_4794;
wire n_4803;
wire n_4802;
wire n_4798;
wire n_5007;
wire n_5006;
wire n_5002;
wire n_5013;
wire n_5014;
wire n_5008;
wire n_4804;
wire n_4877;
wire n_4906;
wire n_4908;
wire n_4904;
wire n_4813;
wire n_4819;
wire n_4909;
wire n_4832;
wire n_4839;
wire n_4915;
wire n_4848;
wire n_4854;
wire n_4922;
wire n_4863;
wire n_4869;
wire n_5016;
wire n_4926;
wire n_4921;
wire n_4919;
wire n_4871;
wire n_4901;
wire n_4880;
wire n_4882;
wire n_4881;
wire n_4941;
wire n_4916;
wire n_4914;
wire n_4912;
wire n_4891;
wire n_4893;
wire n_4887;
wire n_4872;
wire n_4884;
wire n_4878;
wire n_4879;
wire n_4994;
wire n_4883;
wire n_4899;
wire n_4885;
wire n_4961;
wire n_4888;
wire n_4892;
wire n_4895;
wire n_4967;
wire n_4898;
wire n_4932;
wire n_4900;
wire n_4942;
wire n_5096;
wire n_4936;
wire n_4993;
wire n_4902;
wire n_4991;
wire n_4985;
wire n_4903;
wire n_4962;
wire n_4905;
wire n_4907;
wire n_4913;
wire n_4920;
wire n_5015;
wire n_4931;
wire n_4971;
wire n_4999;
wire n_5001;
wire n_4997;
wire n_4935;
wire n_4946;
wire n_4950;
wire n_5029;
wire n_4957;
wire n_5019;
wire n_4966;
wire n_5105;
wire n_5102;
wire n_5101;
wire n_5097;
wire n_5067;
wire n_5076;
wire n_5061;
wire n_4976;
wire n_5030;
wire n_4977;
wire n_5020;
wire n_4981;
wire n_5036;
wire n_4986;
wire n_5047;
wire n_4996;
wire n_5046;
wire n_4998;
wire n_5000;
wire n_5004;
wire n_5005;
wire n_5027;
wire n_5009;
wire n_5012;
wire n_5017;
wire n_5051;
wire n_5042;
wire n_5041;
wire n_5037;
wire n_5086;
wire n_5095;
wire n_5081;
wire n_5026;
wire n_5025;
wire n_5021;
wire n_5022;
wire n_5023;
wire n_5028;
wire n_5034;
wire n_5033;
wire n_5111;
wire n_5035;
wire n_5116;
wire n_5229;
wire n_5115;
wire n_5038;
wire n_5040;
wire n_5142;
wire n_5050;
wire n_5119;
wire n_5139;
wire n_5141;
wire n_5136;
wire n_5056;
wire n_5134;
wire n_5066;
wire n_5071;
wire n_5082;
wire n_5091;
wire n_5234;
wire n_5155;
wire n_5153;
wire n_5149;
wire n_5106;
wire n_5122;
wire n_5123;
wire n_5120;
wire n_5113;
wire n_5146;
wire n_5148;
wire n_5143;
wire n_5117;
wire n_5129;
wire n_5121;
wire n_5126;
wire n_5125;
wire n_5279;
wire n_5236;
wire n_5232;
wire n_5177;
wire n_5172;
wire n_5163;
wire n_5127;
wire n_5128;
wire n_5160;
wire n_5132;
wire n_5182;
wire n_5133;
wire n_5162;
wire n_5135;
wire n_5196;
wire n_5138;
wire n_5140;
wire n_5144;
wire n_5147;
wire n_5181;
wire n_5150;
wire n_5154;
wire n_5207;
wire n_5217;
wire n_5197;
wire n_5227;
wire n_5156;
wire n_5222;
wire n_5218;
wire n_5158;
wire n_5161;
wire n_5283;
wire n_5167;
wire n_5171;
wire n_5272;
wire n_5187;
wire n_5251;
wire n_5192;
wire n_5240;
wire n_5261;
wire n_5264;
wire n_5258;
wire n_5202;
wire n_5212;
wire n_5262;
wire n_5221;
wire n_5243;
wire n_5230;
wire n_5242;
wire n_5233;
wire n_5235;
wire n_5278;
wire n_5276;
wire n_5273;
wire n_5294;
wire n_5245;
wire n_5244;
wire n_5269;
wire n_5271;
wire n_5265;
wire n_5237;
wire n_5249;
wire n_5241;
wire n_5293;
wire n_5248;
wire n_5252;
wire n_5250;
wire n_5253;
wire n_5257;
wire n_5256;
wire n_5255;
wire n_5354;
wire n_5355;
wire n_5350;
wire n_5363;
wire n_5365;
wire n_5360;
wire n_5259;
wire n_5263;
wire n_5313;
wire n_5266;
wire n_5270;
wire n_5274;
wire n_5277;
wire n_5332;
wire n_5328;
wire n_5318;
wire n_5346;
wire n_5317;
wire n_5312;
wire n_5303;
wire n_5359;
wire n_5292;
wire n_5284;
wire n_5282;
wire n_5288;
wire n_5356;
wire n_5298;
wire n_5333;
wire n_5302;
wire n_5349;
wire n_5308;
wire n_5345;
wire n_5323;
wire n_5329;
wire n_5366;
wire n_5344;
wire n_5343;
wire n_5338;
wire n_5340;
wire n_5342;
wire n_5386;
wire n_5347;
wire n_5348;
wire n_5370;
wire n_5376;
wire n_5377;
wire n_5373;
wire n_5352;
wire n_5353;
wire n_5407;
wire n_5361;
wire n_5362;
wire n_5371;
wire n_5449;
wire n_5391;
wire n_5385;
wire n_5381;
wire n_5401;
wire n_5406;
wire n_5396;
wire n_5367;
wire n_5411;
wire n_5369;
wire n_5415;
wire n_5420;
wire n_5417;
wire n_5374;
wire n_5375;
wire n_5380;
wire n_5456;
wire n_5458;
wire n_5452;
wire n_5382;
wire n_5448;
wire n_5397;
wire n_5405;
wire n_5416;
wire n_5472;
wire n_5464;
wire n_5462;
wire n_5460;
wire n_5441;
wire n_5436;
wire n_5431;
wire n_5447;
wire n_5451;
wire n_5443;
wire n_5421;
wire n_5432;
wire n_5435;
wire n_5459;
wire n_5446;
wire n_5450;
wire n_5463;
wire n_5455;
wire n_5457;
wire n_5461;
wire n_5471;
wire n_5469;
wire n_5479;
wire n_5473;
wire n_5476;
wire n_5482;
wire n_5730;
wire n_5484;
wire n_5490;
wire n_5485;
wire n_5734;
wire n_5486;
wire n_5731;
wire n_5729;
wire n_5728;
wire n_5727;
wire n_5725;
wire n_5722;
wire n_5715;
wire n_5711;
wire n_5706;
wire n_5700;
wire n_5696;
wire n_5691;
wire n_5685;
wire n_5680;
wire n_5675;
wire n_5670;
wire n_5667;
wire n_5665;
wire n_5663;
wire n_5659;
wire n_5657;
wire n_5655;
wire n_5652;
wire n_5650;
wire n_5648;
wire n_5645;
wire n_5643;
wire n_5641;
wire n_5639;
wire n_5634;
wire n_5628;
wire n_5624;
wire n_5615;
wire n_5609;
wire n_5604;
wire n_5599;
wire n_5594;
wire n_5588;
wire n_5584;
wire n_5582;
wire n_5578;
wire n_5576;
wire n_5573;
wire n_5571;
wire n_5569;
wire n_5567;
wire n_5564;
wire n_5562;
wire n_5558;
wire n_5556;
wire n_5554;
wire n_5551;
wire n_5549;
wire n_5547;
wire n_5545;
wire n_5542;
wire n_5535;
wire n_5531;
wire n_5525;
wire n_5519;
wire n_5511;
wire n_5505;
wire n_5500;
wire n_5737;
wire n_5735;
wire n_5504;
wire n_5736;
wire n_5510;
wire n_5515;
wire n_5520;
wire n_5530;
wire n_5534;
wire n_5540;
wire n_5544;
wire n_5546;
wire n_5548;
wire n_5550;
wire n_5552;
wire n_5555;
wire n_5557;
wire n_5561;
wire n_5563;
wire n_5565;
wire n_5568;
wire n_5570;
wire n_5572;
wire n_5575;
wire n_5577;
wire n_5579;
wire n_5583;
wire n_5585;
wire n_5589;
wire n_5598;
wire n_5600;
wire n_5608;
wire n_5614;
wire n_5619;
wire n_5625;
wire n_5629;
wire n_5636;
wire n_5640;
wire n_5642;
wire n_5644;
wire n_5646;
wire n_5649;
wire n_5651;
wire n_5654;
wire n_5656;
wire n_5658;
wire n_5662;
wire n_5664;
wire n_5666;
wire n_5669;
wire n_5671;
wire n_5679;
wire n_5681;
wire n_5690;
wire n_5695;
wire n_5699;
wire n_5705;
wire n_5710;
wire n_5714;
wire n_5720;
wire n_5723;
wire n_5726;
wire n_5733;
wire n_5738;
wire n_5741;
wire n_5746;
wire n_5744;
wire n_5749;


INV_X1 i_5047 (.ZN (n_5767), .A (inputB[24]));
INV_X1 i_5046 (.ZN (n_5762), .A (inputB[17]));
INV_X1 i_5045 (.ZN (n_5758), .A (inputB[11]));
INV_X1 i_5043 (.ZN (n_5757), .A (inputB[9]));
INV_X1 i_5042 (.ZN (n_5756), .A (inputB[3]));
INV_X1 i_5041 (.ZN (n_5755), .A (inputB[2]));
INV_X1 i_5039 (.ZN (n_5754), .A (inputB[1]));
INV_X1 i_5038 (.ZN (n_5753), .A (inputA[31]));
INV_X1 i_5037 (.ZN (n_5751), .A (inputA[30]));
INV_X1 i_5035 (.ZN (n_5750), .A (inputA[29]));
NAND2_X1 i_5034 (.ZN (n_5749), .A1 (inputB[29]), .A2 (inputA[31]));
AND2_X1 i_5033 (.ZN (n_5748), .A1 (inputB[30]), .A2 (inputA[30]));
NOR2_X1 i_5031 (.ZN (n_5746), .A1 (n_5749), .A2 (n_5748));
NAND2_X1 i_5030 (.ZN (n_5745), .A1 (inputB[31]), .A2 (inputA[29]));
INV_X1 i_5029 (.ZN (n_5744), .A (n_5745));
AOI21_X1 i_5027 (.ZN (n_5743), .A (n_5746), .B1 (n_5749), .B2 (n_5748));
AOI21_X1 i_5026 (.ZN (n_5742), .A (n_5746), .B1 (n_5744), .B2 (n_5743));
AOI21_X1 i_5025 (.ZN (n_5741), .A (n_127), .B1 (n_126), .B2 (n_5742));
INV_X1 i_5023 (.ZN (n_5738), .A (n_5741));
NAND3_X1 i_5022 (.ZN (n_5737), .A1 (inputB[31]), .A2 (inputA[31]), .A3 (n_5738));
AOI21_X1 i_5021 (.ZN (n_5736), .A (n_5738), .B1 (inputB[31]), .B2 (inputA[31]));
INV_X1 i_5019 (.ZN (n_5735), .A (n_5736));
NAND2_X1 i_5018 (.ZN (n_5734), .A1 (inputB[0]), .A2 (inputA[2]));
AND2_X1 i_5017 (.ZN (result[0]), .A1 (inputB[0]), .A2 (inputA[0]));
NAND2_X1 i_5015 (.ZN (n_5733), .A1 (n_5755), .A2 (result[0]));
NAND2_X1 i_5014 (.ZN (n_5731), .A1 (inputB[1]), .A2 (inputA[1]));
INV_X1 i_5013 (.ZN (n_5730), .A (n_5731));
NAND2_X1 i_5011 (.ZN (n_5729), .A1 (inputB[2]), .A2 (inputA[0]));
AOI22_X1 i_5010 (.ZN (n_5728), .A1 (n_5734), .A2 (n_5733), .B1 (n_5731), .B2 (n_5729));
AOI21_X1 i_5009 (.ZN (n_5727), .A (n_129), .B1 (n_128), .B2 (n_5728));
INV_X1 i_5007 (.ZN (n_5726), .A (n_5727));
AOI21_X1 i_5006 (.ZN (n_5725), .A (n_131), .B1 (n_130), .B2 (n_5726));
INV_X1 i_5005 (.ZN (n_5723), .A (n_5725));
AOI21_X1 i_5003 (.ZN (n_5722), .A (n_133), .B1 (n_132), .B2 (n_5723));
INV_X1 i_5002 (.ZN (n_5720), .A (n_5722));
AOI21_X1 i_5001 (.ZN (n_5715), .A (n_135), .B1 (n_134), .B2 (n_5720));
INV_X1 i_5000 (.ZN (n_5714), .A (n_5715));
AOI21_X1 i_4999 (.ZN (n_5711), .A (n_137), .B1 (n_136), .B2 (n_5714));
INV_X1 i_4998 (.ZN (n_5710), .A (n_5711));
AOI21_X1 i_4997 (.ZN (n_5706), .A (n_139), .B1 (n_138), .B2 (n_5710));
INV_X1 i_4996 (.ZN (n_5705), .A (n_5706));
AOI21_X1 i_4995 (.ZN (n_5700), .A (n_141), .B1 (n_140), .B2 (n_5705));
INV_X1 i_4994 (.ZN (n_5699), .A (n_5700));
AOI21_X1 i_4993 (.ZN (n_5696), .A (n_143), .B1 (n_142), .B2 (n_5699));
INV_X1 i_4992 (.ZN (n_5695), .A (n_5696));
AOI21_X1 i_4991 (.ZN (n_5691), .A (n_145), .B1 (n_144), .B2 (n_5695));
INV_X1 i_4990 (.ZN (n_5690), .A (n_5691));
AOI21_X1 i_4989 (.ZN (n_5685), .A (n_147), .B1 (n_146), .B2 (n_5690));
INV_X1 i_4988 (.ZN (n_5681), .A (n_5685));
AOI21_X1 i_4987 (.ZN (n_5680), .A (n_149), .B1 (n_148), .B2 (n_5681));
INV_X1 i_4986 (.ZN (n_5679), .A (n_5680));
AOI21_X1 i_4985 (.ZN (n_5675), .A (n_151), .B1 (n_150), .B2 (n_5679));
INV_X1 i_4984 (.ZN (n_5671), .A (n_5675));
AOI21_X1 i_4983 (.ZN (n_5670), .A (n_153), .B1 (n_152), .B2 (n_5671));
INV_X1 i_4982 (.ZN (n_5669), .A (n_5670));
AOI21_X1 i_4981 (.ZN (n_5667), .A (n_155), .B1 (n_154), .B2 (n_5669));
INV_X1 i_4980 (.ZN (n_5666), .A (n_5667));
AOI21_X1 i_4979 (.ZN (n_5665), .A (n_157), .B1 (n_156), .B2 (n_5666));
INV_X1 i_4978 (.ZN (n_5664), .A (n_5665));
AOI21_X1 i_4977 (.ZN (n_5663), .A (n_159), .B1 (n_158), .B2 (n_5664));
INV_X1 i_4976 (.ZN (n_5662), .A (n_5663));
AOI21_X1 i_4975 (.ZN (n_5659), .A (n_161), .B1 (n_160), .B2 (n_5662));
INV_X1 i_4974 (.ZN (n_5658), .A (n_5659));
AOI21_X1 i_4973 (.ZN (n_5657), .A (n_163), .B1 (n_162), .B2 (n_5658));
INV_X1 i_4972 (.ZN (n_5656), .A (n_5657));
AOI21_X1 i_4971 (.ZN (n_5655), .A (n_165), .B1 (n_164), .B2 (n_5656));
INV_X1 i_4970 (.ZN (n_5654), .A (n_5655));
AOI21_X1 i_4969 (.ZN (n_5652), .A (n_167), .B1 (n_166), .B2 (n_5654));
INV_X1 i_4968 (.ZN (n_5651), .A (n_5652));
AOI21_X1 i_4967 (.ZN (n_5650), .A (n_169), .B1 (n_168), .B2 (n_5651));
INV_X1 i_4966 (.ZN (n_5649), .A (n_5650));
AOI21_X1 i_4965 (.ZN (n_5648), .A (n_171), .B1 (n_170), .B2 (n_5649));
INV_X1 i_4964 (.ZN (n_5646), .A (n_5648));
AOI21_X1 i_4963 (.ZN (n_5645), .A (n_173), .B1 (n_172), .B2 (n_5646));
INV_X1 i_4962 (.ZN (n_5644), .A (n_5645));
AOI21_X1 i_4961 (.ZN (n_5643), .A (n_175), .B1 (n_174), .B2 (n_5644));
INV_X1 i_4960 (.ZN (n_5642), .A (n_5643));
AOI21_X1 i_4959 (.ZN (n_5641), .A (n_177), .B1 (n_176), .B2 (n_5642));
INV_X1 i_4958 (.ZN (n_5640), .A (n_5641));
AOI21_X1 i_4957 (.ZN (n_5639), .A (n_179), .B1 (n_178), .B2 (n_5640));
INV_X1 i_4955 (.ZN (n_5636), .A (n_5639));
AOI21_X1 i_4954 (.ZN (n_5634), .A (n_181), .B1 (n_180), .B2 (n_5636));
INV_X1 i_4953 (.ZN (n_5629), .A (n_5634));
AOI21_X1 i_4951 (.ZN (n_5628), .A (n_183), .B1 (n_182), .B2 (n_5629));
INV_X1 i_4950 (.ZN (n_5625), .A (n_5628));
AOI21_X1 i_4949 (.ZN (n_5624), .A (n_185), .B1 (n_184), .B2 (n_5625));
INV_X1 i_4947 (.ZN (n_5619), .A (n_5624));
AOI21_X1 i_4946 (.ZN (n_5615), .A (n_187), .B1 (n_186), .B2 (n_5619));
INV_X1 i_4945 (.ZN (n_5614), .A (n_5615));
AOI21_X1 i_4943 (.ZN (n_5609), .A (n_189), .B1 (n_188), .B2 (n_5614));
INV_X1 i_4942 (.ZN (n_5608), .A (n_5609));
AOI21_X1 i_4941 (.ZN (n_5604), .A (n_191), .B1 (n_190), .B2 (n_5608));
INV_X1 i_4939 (.ZN (n_5600), .A (n_5604));
AOI21_X1 i_4938 (.ZN (n_5599), .A (n_193), .B1 (n_192), .B2 (n_5600));
INV_X1 i_4937 (.ZN (n_5598), .A (n_5599));
AOI21_X1 i_4935 (.ZN (n_5594), .A (n_195), .B1 (n_194), .B2 (n_5598));
INV_X1 i_4934 (.ZN (n_5589), .A (n_5594));
AOI21_X1 i_4933 (.ZN (n_5588), .A (n_197), .B1 (n_196), .B2 (n_5589));
INV_X1 i_4931 (.ZN (n_5585), .A (n_5588));
AOI21_X1 i_4930 (.ZN (n_5584), .A (n_199), .B1 (n_198), .B2 (n_5585));
INV_X1 i_4929 (.ZN (n_5583), .A (n_5584));
AOI21_X1 i_4927 (.ZN (n_5582), .A (n_201), .B1 (n_200), .B2 (n_5583));
INV_X1 i_4926 (.ZN (n_5579), .A (n_5582));
AOI21_X1 i_4925 (.ZN (n_5578), .A (n_203), .B1 (n_202), .B2 (n_5579));
INV_X1 i_4923 (.ZN (n_5577), .A (n_5578));
AOI21_X1 i_4922 (.ZN (n_5576), .A (n_205), .B1 (n_204), .B2 (n_5577));
INV_X1 i_4921 (.ZN (n_5575), .A (n_5576));
AOI21_X1 i_4919 (.ZN (n_5573), .A (n_207), .B1 (n_206), .B2 (n_5575));
INV_X1 i_4918 (.ZN (n_5572), .A (n_5573));
AOI21_X1 i_4917 (.ZN (n_5571), .A (n_209), .B1 (n_208), .B2 (n_5572));
INV_X1 i_4915 (.ZN (n_5570), .A (n_5571));
AOI21_X1 i_4914 (.ZN (n_5569), .A (n_211), .B1 (n_210), .B2 (n_5570));
INV_X1 i_4913 (.ZN (n_5568), .A (n_5569));
AOI21_X1 i_4911 (.ZN (n_5567), .A (n_213), .B1 (n_212), .B2 (n_5568));
INV_X1 i_4910 (.ZN (n_5565), .A (n_5567));
AOI21_X1 i_4909 (.ZN (n_5564), .A (n_215), .B1 (n_214), .B2 (n_5565));
INV_X1 i_4908 (.ZN (n_5563), .A (n_5564));
AOI21_X1 i_4907 (.ZN (n_5562), .A (n_217), .B1 (n_216), .B2 (n_5563));
INV_X1 i_4906 (.ZN (n_5561), .A (n_5562));
AOI21_X1 i_4905 (.ZN (n_5558), .A (n_219), .B1 (n_218), .B2 (n_5561));
INV_X1 i_4904 (.ZN (n_5557), .A (n_5558));
AOI21_X1 i_4903 (.ZN (n_5556), .A (n_221), .B1 (n_220), .B2 (n_5557));
INV_X1 i_4902 (.ZN (n_5555), .A (n_5556));
AOI21_X1 i_4901 (.ZN (n_5554), .A (n_223), .B1 (n_222), .B2 (n_5555));
INV_X1 i_4900 (.ZN (n_5552), .A (n_5554));
AOI21_X1 i_4899 (.ZN (n_5551), .A (n_225), .B1 (n_224), .B2 (n_5552));
INV_X1 i_4898 (.ZN (n_5550), .A (n_5551));
AOI21_X1 i_4897 (.ZN (n_5549), .A (n_227), .B1 (n_226), .B2 (n_5550));
INV_X1 i_4896 (.ZN (n_5548), .A (n_5549));
AOI21_X1 i_4895 (.ZN (n_5547), .A (n_229), .B1 (n_228), .B2 (n_5548));
INV_X1 i_4894 (.ZN (n_5546), .A (n_5547));
AOI21_X1 i_4893 (.ZN (n_5545), .A (n_231), .B1 (n_230), .B2 (n_5546));
INV_X1 i_4892 (.ZN (n_5544), .A (n_5545));
AOI21_X1 i_4891 (.ZN (n_5542), .A (n_233), .B1 (n_232), .B2 (n_5544));
INV_X1 i_4890 (.ZN (n_5540), .A (n_5542));
AOI21_X1 i_4889 (.ZN (n_5535), .A (n_235), .B1 (n_234), .B2 (n_5540));
INV_X1 i_4888 (.ZN (n_5534), .A (n_5535));
AOI21_X1 i_4887 (.ZN (n_5531), .A (n_237), .B1 (n_236), .B2 (n_5534));
INV_X1 i_4886 (.ZN (n_5530), .A (n_5531));
AOI21_X1 i_4885 (.ZN (n_5525), .A (n_239), .B1 (n_238), .B2 (n_5530));
INV_X1 i_4884 (.ZN (n_5520), .A (n_5525));
AOI21_X1 i_4883 (.ZN (n_5519), .A (n_241), .B1 (n_240), .B2 (n_5520));
INV_X1 i_4882 (.ZN (n_5515), .A (n_5519));
AOI21_X1 i_4881 (.ZN (n_5511), .A (n_243), .B1 (n_242), .B2 (n_5515));
INV_X1 i_4880 (.ZN (n_5510), .A (n_5511));
AOI21_X1 i_4879 (.ZN (n_5505), .A (n_245), .B1 (n_244), .B2 (n_5510));
AOI21_X1 i_4878 (.ZN (n_5504), .A (n_5736), .B1 (n_5737), .B2 (n_5505));
INV_X1 i_4877 (.ZN (result[63]), .A (n_5504));
NAND2_X1 i_4876 (.ZN (n_5500), .A1 (n_5737), .A2 (n_5735));
XOR2_X1 i_4875 (.Z (result[62]), .A (n_5505), .B (n_5500));
XNOR2_X1 i_4874 (.ZN (result[61]), .A (n_244), .B (n_5511));
XNOR2_X1 i_4873 (.ZN (result[60]), .A (n_242), .B (n_5519));
XNOR2_X1 i_4872 (.ZN (result[59]), .A (n_240), .B (n_5525));
XNOR2_X1 i_4871 (.ZN (result[58]), .A (n_238), .B (n_5531));
XNOR2_X1 i_4870 (.ZN (result[57]), .A (n_236), .B (n_5535));
XNOR2_X1 i_4869 (.ZN (result[56]), .A (n_234), .B (n_5542));
XNOR2_X1 i_4868 (.ZN (result[55]), .A (n_232), .B (n_5545));
XNOR2_X1 i_4867 (.ZN (result[54]), .A (n_230), .B (n_5547));
XNOR2_X1 i_4866 (.ZN (result[53]), .A (n_228), .B (n_5549));
XNOR2_X1 i_4864 (.ZN (result[52]), .A (n_226), .B (n_5551));
XNOR2_X1 i_4863 (.ZN (result[51]), .A (n_224), .B (n_5554));
XNOR2_X1 i_4862 (.ZN (result[50]), .A (n_222), .B (n_5556));
XNOR2_X1 i_4860 (.ZN (result[49]), .A (n_220), .B (n_5558));
XNOR2_X1 i_4859 (.ZN (result[48]), .A (n_218), .B (n_5562));
XNOR2_X1 i_4858 (.ZN (result[47]), .A (n_216), .B (n_5564));
XNOR2_X1 i_4856 (.ZN (result[46]), .A (n_214), .B (n_5567));
XNOR2_X1 i_4855 (.ZN (result[45]), .A (n_212), .B (n_5569));
XNOR2_X1 i_4854 (.ZN (result[44]), .A (n_210), .B (n_5571));
XNOR2_X1 i_4852 (.ZN (result[43]), .A (n_208), .B (n_5573));
XNOR2_X1 i_4851 (.ZN (result[42]), .A (n_206), .B (n_5576));
XNOR2_X1 i_4850 (.ZN (result[41]), .A (n_204), .B (n_5578));
XNOR2_X1 i_4848 (.ZN (result[40]), .A (n_202), .B (n_5582));
XNOR2_X1 i_4847 (.ZN (result[39]), .A (n_200), .B (n_5584));
XNOR2_X1 i_4846 (.ZN (result[38]), .A (n_198), .B (n_5588));
XNOR2_X1 i_4844 (.ZN (result[37]), .A (n_196), .B (n_5594));
XNOR2_X1 i_4843 (.ZN (result[36]), .A (n_194), .B (n_5599));
XNOR2_X1 i_4842 (.ZN (result[35]), .A (n_192), .B (n_5604));
XNOR2_X1 i_4840 (.ZN (result[34]), .A (n_190), .B (n_5609));
XNOR2_X1 i_4839 (.ZN (result[33]), .A (n_188), .B (n_5615));
XNOR2_X1 i_4838 (.ZN (result[32]), .A (n_186), .B (n_5624));
XNOR2_X1 i_4836 (.ZN (result[31]), .A (n_184), .B (n_5628));
XNOR2_X1 i_4835 (.ZN (result[30]), .A (n_182), .B (n_5634));
XNOR2_X1 i_4834 (.ZN (result[29]), .A (n_180), .B (n_5639));
XNOR2_X1 i_4832 (.ZN (result[28]), .A (n_178), .B (n_5641));
XNOR2_X1 i_4831 (.ZN (result[27]), .A (n_176), .B (n_5643));
XNOR2_X1 i_4830 (.ZN (result[26]), .A (n_174), .B (n_5645));
XNOR2_X1 i_4828 (.ZN (result[25]), .A (n_172), .B (n_5648));
XNOR2_X1 i_4827 (.ZN (result[24]), .A (n_170), .B (n_5650));
XNOR2_X1 i_4826 (.ZN (result[23]), .A (n_168), .B (n_5652));
XNOR2_X1 i_4824 (.ZN (result[22]), .A (n_166), .B (n_5655));
XNOR2_X1 i_4823 (.ZN (result[21]), .A (n_164), .B (n_5657));
XNOR2_X1 i_4822 (.ZN (result[20]), .A (n_162), .B (n_5659));
XNOR2_X1 i_4820 (.ZN (result[19]), .A (n_160), .B (n_5663));
XNOR2_X1 i_4819 (.ZN (result[18]), .A (n_158), .B (n_5665));
XNOR2_X1 i_4818 (.ZN (result[17]), .A (n_156), .B (n_5667));
XNOR2_X1 i_4817 (.ZN (result[16]), .A (n_154), .B (n_5670));
XNOR2_X1 i_4816 (.ZN (result[15]), .A (n_152), .B (n_5675));
XNOR2_X1 i_4815 (.ZN (result[14]), .A (n_150), .B (n_5680));
XNOR2_X1 i_4814 (.ZN (result[13]), .A (n_148), .B (n_5685));
XNOR2_X1 i_4813 (.ZN (result[12]), .A (n_146), .B (n_5691));
XNOR2_X1 i_4812 (.ZN (result[11]), .A (n_144), .B (n_5696));
XNOR2_X1 i_4811 (.ZN (result[10]), .A (n_142), .B (n_5700));
XNOR2_X1 i_4810 (.ZN (result[9]), .A (n_140), .B (n_5706));
XNOR2_X1 i_4809 (.ZN (result[8]), .A (n_138), .B (n_5711));
XNOR2_X1 i_4808 (.ZN (result[7]), .A (n_136), .B (n_5715));
XNOR2_X1 i_4807 (.ZN (result[6]), .A (n_134), .B (n_5722));
XNOR2_X1 i_4806 (.ZN (result[5]), .A (n_132), .B (n_5725));
XNOR2_X1 i_4805 (.ZN (result[4]), .A (n_130), .B (n_5727));
XOR2_X1 i_4804 (.Z (result[3]), .A (n_128), .B (n_5728));
NOR2_X1 i_4803 (.ZN (n_5496), .A1 (n_5731), .A2 (n_5729));
INV_X1 i_4802 (.ZN (n_5495), .A (n_5496));
AOI21_X1 i_4801 (.ZN (n_5490), .A (n_5496), .B1 (n_5731), .B2 (n_5729));
NAND2_X1 i_4800 (.ZN (n_5486), .A1 (result[0]), .A2 (n_5730));
XOR2_X1 i_4799 (.Z (n_5485), .A (n_5734), .B (n_5486));
XOR2_X1 i_4798 (.Z (result[2]), .A (n_5490), .B (n_5485));
AOI22_X1 i_4797 (.ZN (n_5484), .A1 (inputB[1]), .A2 (inputA[0]), .B1 (inputB[0]), .B2 (inputA[1]));
AOI21_X1 i_4796 (.ZN (result[1]), .A (n_5484), .B1 (result[0]), .B2 (n_5730));
NAND3_X1 i_4795 (.ZN (n_5483), .A1 (inputB[2]), .A2 (inputA[2]), .A3 (n_5730));
AOI22_X1 i_4794 (.ZN (n_5482), .A1 (inputB[2]), .A2 (inputA[1]), .B1 (inputB[1]), .B2 (inputA[2]));
INV_X1 i_4793 (.ZN (n_5481), .A (n_5482));
NAND2_X1 i_4792 (.ZN (n_5480), .A1 (inputB[3]), .A2 (inputA[0]));
AOI21_X1 i_4791 (.ZN (n_1030), .A (n_5482), .B1 (n_5483), .B2 (n_5480));
AOI22_X1 i_4790 (.ZN (n_5479), .A1 (inputB[1]), .A2 (inputA[3]), .B1 (inputB[0]), .B2 (inputA[4]));
NAND2_X1 i_4789 (.ZN (n_5478), .A1 (inputB[0]), .A2 (inputA[3]));
INV_X1 i_4788 (.ZN (n_5477), .A (n_5478));
AOI21_X1 i_4787 (.ZN (n_5476), .A (n_5496), .B1 (inputB[1]), .B2 (inputA[4]));
NOR2_X1 i_4786 (.ZN (n_1046), .A1 (n_5478), .A2 (n_5476));
NAND2_X1 i_4785 (.ZN (n_5473), .A1 (inputA[4]), .A2 (n_5477));
OAI22_X1 i_4784 (.ZN (n_1045), .A1 (n_5479), .A2 (n_1046), .B1 (n_5495), .B2 (n_5473));
NAND2_X1 i_4783 (.ZN (n_5472), .A1 (inputB[3]), .A2 (inputA[2]));
INV_X1 i_4782 (.ZN (n_5471), .A (n_5472));
NAND3_X1 i_4781 (.ZN (n_5470), .A1 (inputB[2]), .A2 (inputA[1]), .A3 (n_5471));
AOI22_X1 i_4780 (.ZN (n_5469), .A1 (inputB[2]), .A2 (inputA[2]), .B1 (inputB[3]), .B2 (inputA[1]));
INV_X1 i_4779 (.ZN (n_5466), .A (n_5469));
NAND2_X1 i_4778 (.ZN (n_5465), .A1 (inputB[4]), .A2 (inputA[0]));
AOI21_X1 i_4777 (.ZN (n_1040), .A (n_5469), .B1 (n_5470), .B2 (n_5465));
NAND2_X1 i_4776 (.ZN (n_5464), .A1 (inputB[4]), .A2 (inputA[1]));
INV_X1 i_4775 (.ZN (n_5463), .A (n_5464));
NAND2_X1 i_4774 (.ZN (n_5462), .A1 (n_5471), .A2 (n_5463));
OAI21_X1 i_4773 (.ZN (n_5461), .A (n_5462), .B1 (n_5471), .B2 (n_5463));
NAND2_X1 i_4772 (.ZN (n_5460), .A1 (inputB[5]), .A2 (inputA[0]));
XOR2_X1 i_4771 (.Z (n_1056), .A (n_5461), .B (n_5460));
AND2_X1 i_4770 (.ZN (n_5459), .A1 (inputB[1]), .A2 (inputA[5]));
AOI21_X1 i_4769 (.ZN (n_5458), .A (n_5459), .B1 (inputB[2]), .B2 (inputA[4]));
INV_X1 i_4768 (.ZN (n_5457), .A (n_5458));
NAND3_X1 i_4767 (.ZN (n_5456), .A1 (inputB[2]), .A2 (inputA[4]), .A3 (n_5459));
NAND2_X1 i_4765 (.ZN (n_5455), .A1 (n_5457), .A2 (n_5456));
NAND2_X1 i_4764 (.ZN (n_5452), .A1 (inputB[3]), .A2 (inputA[3]));
XOR2_X1 i_4763 (.Z (n_1084), .A (n_5455), .B (n_5452));
AOI22_X1 i_4761 (.ZN (n_5451), .A1 (inputB[4]), .A2 (inputA[2]), .B1 (inputB[5]), .B2 (inputA[1]));
INV_X1 i_4760 (.ZN (n_5450), .A (n_5451));
NAND2_X1 i_4759 (.ZN (n_5449), .A1 (inputB[5]), .A2 (inputA[2]));
INV_X1 i_4757 (.ZN (n_5448), .A (n_5449));
NAND2_X1 i_4756 (.ZN (n_5447), .A1 (n_5463), .A2 (n_5448));
NAND2_X1 i_4755 (.ZN (n_5446), .A1 (n_5450), .A2 (n_5447));
NAND2_X1 i_4753 (.ZN (n_5443), .A1 (inputB[6]), .A2 (inputA[0]));
XOR2_X1 i_4752 (.Z (n_1077), .A (n_5446), .B (n_5443));
NAND3_X1 i_4751 (.ZN (n_5441), .A1 (inputB[0]), .A2 (inputA[4]), .A3 (n_5459));
AOI22_X1 i_4749 (.ZN (n_5436), .A1 (inputB[1]), .A2 (inputA[4]), .B1 (inputB[0]), .B2 (inputA[5]));
INV_X1 i_4748 (.ZN (n_5435), .A (n_5436));
NAND2_X1 i_4747 (.ZN (n_5432), .A1 (n_5441), .A2 (n_5435));
NAND2_X1 i_4745 (.ZN (n_5431), .A1 (inputB[2]), .A2 (inputA[3]));
XOR2_X1 i_4744 (.Z (n_5426), .A (n_5432), .B (n_5431));
AOI21_X1 i_4743 (.ZN (n_5421), .A (n_1069), .B1 (n_1068), .B2 (n_5426));
INV_X1 i_4741 (.ZN (n_1072), .A (n_5421));
OAI21_X1 i_4740 (.ZN (n_1078), .A (n_5447), .B1 (n_5451), .B2 (n_5443));
OAI21_X1 i_4739 (.ZN (n_5420), .A (n_5441), .B1 (n_5436), .B2 (n_5431));
AOI22_X1 i_4737 (.ZN (n_5417), .A1 (n_5472), .A2 (n_5464), .B1 (n_5462), .B2 (n_5460));
NOR2_X1 i_4736 (.ZN (n_5416), .A1 (n_5420), .A2 (n_5417));
NAND2_X1 i_4735 (.ZN (n_5415), .A1 (n_5420), .A2 (n_5417));
NAND2_X1 i_4733 (.ZN (n_5411), .A1 (inputB[0]), .A2 (inputA[6]));
OAI21_X1 i_4732 (.ZN (n_1092), .A (n_5415), .B1 (n_5416), .B2 (n_5411));
AND2_X1 i_4731 (.ZN (n_5407), .A1 (inputB[3]), .A2 (inputA[4]));
AOI21_X1 i_4729 (.ZN (n_5406), .A (n_5407), .B1 (inputB[2]), .B2 (inputA[5]));
INV_X1 i_4728 (.ZN (n_5405), .A (n_5406));
NAND3_X1 i_4727 (.ZN (n_5401), .A1 (inputB[2]), .A2 (inputA[5]), .A3 (n_5407));
NAND2_X1 i_4725 (.ZN (n_5397), .A1 (n_5405), .A2 (n_5401));
NAND2_X1 i_4724 (.ZN (n_5396), .A1 (inputB[4]), .A2 (inputA[3]));
XOR2_X1 i_4723 (.Z (n_1113), .A (n_5397), .B (n_5396));
NAND2_X1 i_4721 (.ZN (n_5391), .A1 (inputB[6]), .A2 (inputA[1]));
INV_X1 i_4720 (.ZN (n_5386), .A (n_5391));
NAND2_X1 i_4719 (.ZN (n_5385), .A1 (n_5448), .A2 (n_5386));
OAI21_X1 i_4717 (.ZN (n_5382), .A (n_5385), .B1 (n_5448), .B2 (n_5386));
NAND2_X1 i_4716 (.ZN (n_5381), .A1 (inputB[7]), .A2 (inputA[0]));
XOR2_X1 i_4715 (.Z (n_1106), .A (n_5382), .B (n_5381));
OAI21_X1 i_4714 (.ZN (n_5380), .A (n_5456), .B1 (n_5458), .B2 (n_5452));
AOI21_X1 i_4713 (.ZN (n_5377), .A (n_5380), .B1 (inputB[1]), .B2 (inputA[6]));
NAND3_X1 i_4712 (.ZN (n_5376), .A1 (inputB[1]), .A2 (inputA[6]), .A3 (n_5380));
INV_X1 i_4711 (.ZN (n_5375), .A (n_5376));
NOR2_X1 i_4710 (.ZN (n_5374), .A1 (n_5377), .A2 (n_5375));
NAND2_X1 i_4709 (.ZN (n_5373), .A1 (inputB[0]), .A2 (inputA[7]));
INV_X1 i_4708 (.ZN (n_5371), .A (n_5373));
XOR2_X1 i_4707 (.Z (n_5370), .A (n_5374), .B (n_5371));
XOR2_X1 i_4706 (.Z (n_1128), .A (n_1126), .B (n_5370));
OAI21_X1 i_4705 (.ZN (n_5369), .A (n_5415), .B1 (n_5420), .B2 (n_5417));
XOR2_X1 i_4704 (.Z (n_5368), .A (n_5411), .B (n_5369));
AOI21_X1 i_4703 (.ZN (n_5367), .A (n_1098), .B1 (n_1097), .B2 (n_5368));
INV_X1 i_4702 (.ZN (n_1101), .A (n_5367));
OAI21_X1 i_4701 (.ZN (n_1114), .A (n_5401), .B1 (n_5406), .B2 (n_5396));
AOI22_X1 i_4700 (.ZN (n_1107), .A1 (n_5449), .A2 (n_5391), .B1 (n_5385), .B2 (n_5381));
AND2_X1 i_4699 (.ZN (n_5366), .A1 (inputB[1]), .A2 (inputA[8]));
NAND2_X1 i_4698 (.ZN (n_5365), .A1 (n_5371), .A2 (n_5366));
AOI22_X1 i_4697 (.ZN (n_5363), .A1 (inputB[0]), .A2 (inputA[8]), .B1 (inputB[1]), .B2 (inputA[7]));
INV_X1 i_4696 (.ZN (n_5362), .A (n_5363));
NAND2_X1 i_4695 (.ZN (n_5361), .A1 (n_5365), .A2 (n_5362));
NAND2_X1 i_4694 (.ZN (n_5360), .A1 (inputB[2]), .A2 (inputA[6]));
XOR2_X1 i_4693 (.Z (n_1154), .A (n_5361), .B (n_5360));
NAND2_X1 i_4692 (.ZN (n_5359), .A1 (inputB[4]), .A2 (inputA[5]));
INV_X1 i_4691 (.ZN (n_5356), .A (n_5359));
NAND2_X1 i_4690 (.ZN (n_5355), .A1 (n_5407), .A2 (n_5356));
AOI22_X1 i_4689 (.ZN (n_5354), .A1 (inputB[3]), .A2 (inputA[5]), .B1 (inputB[4]), .B2 (inputA[4]));
INV_X1 i_4688 (.ZN (n_5353), .A (n_5354));
NAND2_X1 i_4687 (.ZN (n_5352), .A1 (n_5355), .A2 (n_5353));
NAND2_X1 i_4686 (.ZN (n_5350), .A1 (inputB[5]), .A2 (inputA[3]));
XOR2_X1 i_4685 (.Z (n_1147), .A (n_5352), .B (n_5350));
OAI21_X1 i_4684 (.ZN (n_5349), .A (n_5376), .B1 (n_5377), .B2 (n_5373));
XOR2_X1 i_4683 (.Z (n_1161), .A (n_1159), .B (n_5349));
AOI21_X1 i_4682 (.ZN (n_5348), .A (n_1127), .B1 (n_1126), .B2 (n_5370));
INV_X1 i_4681 (.ZN (n_1130), .A (n_5348));
AOI21_X1 i_4680 (.ZN (n_5347), .A (n_1132), .B1 (n_1103), .B2 (n_1131));
INV_X1 i_4679 (.ZN (n_1135), .A (n_5347));
NAND2_X1 i_4678 (.ZN (n_5346), .A1 (inputB[7]), .A2 (inputA[2]));
INV_X1 i_4677 (.ZN (n_5345), .A (n_5346));
NAND2_X1 i_4676 (.ZN (n_5344), .A1 (n_5386), .A2 (n_5345));
AOI22_X1 i_4675 (.ZN (n_5343), .A1 (inputB[6]), .A2 (inputA[2]), .B1 (inputB[7]), .B2 (inputA[1]));
INV_X1 i_4674 (.ZN (n_5342), .A (n_5343));
NAND2_X1 i_4673 (.ZN (n_5340), .A1 (n_5344), .A2 (n_5342));
NAND2_X1 i_4672 (.ZN (n_5338), .A1 (inputB[8]), .A2 (inputA[0]));
XOR2_X1 i_4671 (.Z (n_5333), .A (n_5340), .B (n_5338));
XOR2_X1 i_4670 (.Z (n_1166), .A (n_1164), .B (n_5333));
OAI21_X1 i_4669 (.ZN (n_1141), .A (n_5344), .B1 (n_5343), .B2 (n_5338));
AND3_X1 i_4668 (.ZN (n_5332), .A1 (inputB[2]), .A2 (inputA[7]), .A3 (n_5366));
AOI21_X1 i_4667 (.ZN (n_5329), .A (n_5366), .B1 (inputB[2]), .B2 (inputA[7]));
INV_X1 i_4666 (.ZN (n_5328), .A (n_5329));
NOR2_X1 i_4665 (.ZN (n_5323), .A1 (n_5332), .A2 (n_5329));
AND2_X1 i_4664 (.ZN (n_5318), .A1 (inputB[3]), .A2 (inputA[6]));
XOR2_X1 i_4662 (.Z (n_1192), .A (n_5323), .B (n_5318));
NAND2_X1 i_4661 (.ZN (n_5317), .A1 (inputB[8]), .A2 (inputA[1]));
INV_X1 i_4660 (.ZN (n_5313), .A (n_5317));
NAND2_X1 i_4658 (.ZN (n_5312), .A1 (n_5345), .A2 (n_5313));
OAI21_X1 i_4657 (.ZN (n_5308), .A (n_5312), .B1 (n_5345), .B2 (n_5313));
NAND2_X1 i_4656 (.ZN (n_5303), .A1 (inputB[9]), .A2 (inputA[0]));
XOR2_X1 i_4654 (.Z (n_1178), .A (n_5308), .B (n_5303));
AOI21_X1 i_4653 (.ZN (n_5302), .A (n_1160), .B1 (n_1159), .B2 (n_5349));
INV_X1 i_4652 (.ZN (n_1163), .A (n_5302));
AOI21_X1 i_4650 (.ZN (n_5298), .A (n_1165), .B1 (n_1164), .B2 (n_5333));
INV_X1 i_4649 (.ZN (n_1168), .A (n_5298));
NAND2_X1 i_4648 (.ZN (n_5294), .A1 (inputB[5]), .A2 (inputA[4]));
INV_X1 i_4646 (.ZN (n_5293), .A (n_5294));
NAND2_X1 i_4645 (.ZN (n_5292), .A1 (n_5356), .A2 (n_5293));
OAI21_X1 i_4644 (.ZN (n_5288), .A (n_5292), .B1 (n_5356), .B2 (n_5293));
NAND2_X1 i_4642 (.ZN (n_5284), .A1 (inputB[6]), .A2 (inputA[3]));
XOR2_X1 i_4641 (.Z (n_5283), .A (n_5288), .B (n_5284));
XOR2_X1 i_4640 (.Z (n_1207), .A (n_1205), .B (n_5283));
AOI21_X1 i_4638 (.ZN (n_5282), .A (n_1170), .B1 (n_1137), .B2 (n_1169));
INV_X1 i_4637 (.ZN (n_1173), .A (n_5282));
AOI22_X1 i_4636 (.ZN (n_1186), .A1 (n_5359), .A2 (n_5294), .B1 (n_5292), .B2 (n_5284));
AOI22_X1 i_4634 (.ZN (n_1179), .A1 (n_5346), .A2 (n_5317), .B1 (n_5312), .B2 (n_5303));
NAND2_X1 i_4633 (.ZN (n_5279), .A1 (inputB[0]), .A2 (inputA[10]));
AOI21_X1 i_4632 (.ZN (n_5278), .A (n_5332), .B1 (n_5328), .B2 (n_5318));
NAND2_X1 i_4630 (.ZN (n_5277), .A1 (n_5279), .A2 (n_5278));
INV_X1 i_4629 (.ZN (n_5276), .A (n_5277));
OAI21_X1 i_4628 (.ZN (n_5274), .A (n_5277), .B1 (n_5279), .B2 (n_5278));
NAND2_X1 i_4626 (.ZN (n_5273), .A1 (inputB[1]), .A2 (inputA[9]));
XOR2_X1 i_4625 (.Z (n_1244), .A (n_5274), .B (n_5273));
AND2_X1 i_4624 (.ZN (n_5272), .A1 (inputB[3]), .A2 (inputA[7]));
AOI21_X1 i_4622 (.ZN (n_5271), .A (n_5272), .B1 (inputB[2]), .B2 (inputA[8]));
INV_X1 i_4621 (.ZN (n_5270), .A (n_5271));
NAND3_X1 i_4620 (.ZN (n_5269), .A1 (inputB[2]), .A2 (inputA[8]), .A3 (n_5272));
NAND2_X1 i_4618 (.ZN (n_5266), .A1 (n_5270), .A2 (n_5269));
NAND2_X1 i_4617 (.ZN (n_5265), .A1 (inputB[4]), .A2 (inputA[6]));
XOR2_X1 i_4616 (.Z (n_1238), .A (n_5266), .B (n_5265));
AOI22_X1 i_4614 (.ZN (n_5264), .A1 (inputB[8]), .A2 (inputA[2]), .B1 (inputB[9]), .B2 (inputA[1]));
INV_X1 i_4613 (.ZN (n_5263), .A (n_5264));
AND2_X1 i_4612 (.ZN (n_5262), .A1 (inputB[9]), .A2 (inputA[2]));
NAND2_X1 i_4610 (.ZN (n_5261), .A1 (n_5313), .A2 (n_5262));
NAND2_X1 i_4609 (.ZN (n_5259), .A1 (n_5263), .A2 (n_5261));
NAND2_X1 i_4608 (.ZN (n_5258), .A1 (inputB[10]), .A2 (inputA[0]));
XOR2_X1 i_4607 (.Z (n_1224), .A (n_5259), .B (n_5258));
AOI21_X1 i_4606 (.ZN (n_5257), .A (n_5363), .B1 (n_5365), .B2 (n_5360));
AOI21_X1 i_4605 (.ZN (n_5256), .A (n_5354), .B1 (n_5355), .B2 (n_5350));
NOR2_X1 i_4604 (.ZN (n_5255), .A1 (n_5257), .A2 (n_5256));
NAND2_X1 i_4603 (.ZN (n_5253), .A1 (n_5257), .A2 (n_5256));
NAND2_X1 i_4602 (.ZN (n_5252), .A1 (inputB[0]), .A2 (inputA[9]));
OAI21_X1 i_4601 (.ZN (n_5251), .A (n_5253), .B1 (n_5255), .B2 (n_5252));
XOR2_X1 i_4600 (.Z (n_1253), .A (n_1251), .B (n_5251));
OAI21_X1 i_4599 (.ZN (n_5250), .A (n_5253), .B1 (n_5257), .B2 (n_5256));
XOR2_X1 i_4598 (.Z (n_5249), .A (n_5252), .B (n_5250));
AOI21_X1 i_4597 (.ZN (n_5248), .A (n_1211), .B1 (n_1210), .B2 (n_5249));
INV_X1 i_4596 (.ZN (n_1214), .A (n_5248));
NAND2_X1 i_4595 (.ZN (n_5245), .A1 (inputB[7]), .A2 (inputA[3]));
AOI22_X1 i_4594 (.ZN (n_5244), .A1 (inputB[5]), .A2 (inputA[5]), .B1 (inputB[6]), .B2 (inputA[4]));
NAND2_X1 i_4593 (.ZN (n_5243), .A1 (inputB[6]), .A2 (inputA[5]));
INV_X1 i_4592 (.ZN (n_5242), .A (n_5243));
AOI21_X1 i_4591 (.ZN (n_5241), .A (n_5244), .B1 (n_5293), .B2 (n_5242));
XNOR2_X1 i_4590 (.ZN (n_5240), .A (n_5245), .B (n_5241));
XOR2_X1 i_4589 (.Z (n_1258), .A (n_1256), .B (n_5240));
XOR2_X1 i_4588 (.Z (n_5238), .A (n_1210), .B (n_5249));
AOI21_X1 i_4587 (.ZN (n_5237), .A (n_1216), .B1 (n_1215), .B2 (n_5238));
INV_X1 i_4586 (.ZN (n_1219), .A (n_5237));
OAI21_X1 i_4585 (.ZN (n_1239), .A (n_5269), .B1 (n_5271), .B2 (n_5265));
OAI22_X1 i_4584 (.ZN (n_1232), .A1 (n_5294), .A2 (n_5243), .B1 (n_5245), .B2 (n_5244));
OAI22_X1 i_4583 (.ZN (n_1245), .A1 (n_5279), .A2 (n_5278), .B1 (n_5276), .B2 (n_5273));
AOI22_X1 i_4582 (.ZN (n_5236), .A1 (inputB[0]), .A2 (inputA[11]), .B1 (inputB[1]), .B2 (inputA[10]));
INV_X1 i_4581 (.ZN (n_5235), .A (n_5236));
NAND2_X1 i_4580 (.ZN (n_5234), .A1 (inputB[1]), .A2 (inputA[11]));
OAI21_X1 i_4579 (.ZN (n_5233), .A (n_5235), .B1 (n_5279), .B2 (n_5234));
NAND2_X1 i_4578 (.ZN (n_5232), .A1 (inputB[2]), .A2 (inputA[9]));
XOR2_X1 i_4577 (.Z (n_1296), .A (n_5233), .B (n_5232));
NAND2_X1 i_4576 (.ZN (n_5230), .A1 (inputB[7]), .A2 (inputA[4]));
INV_X1 i_4575 (.ZN (n_5229), .A (n_5230));
NAND2_X1 i_4574 (.ZN (n_5227), .A1 (n_5242), .A2 (n_5229));
NAND2_X1 i_4573 (.ZN (n_5222), .A1 (n_5243), .A2 (n_5230));
AND2_X1 i_4572 (.ZN (n_5221), .A1 (n_5227), .A2 (n_5222));
AND2_X1 i_4571 (.ZN (n_5218), .A1 (inputB[8]), .A2 (inputA[3]));
XOR2_X1 i_4570 (.Z (n_1282), .A (n_5221), .B (n_5218));
AOI21_X1 i_4569 (.ZN (n_5217), .A (n_5262), .B1 (inputB[10]), .B2 (inputA[1]));
INV_X1 i_4568 (.ZN (n_5212), .A (n_5217));
NAND3_X1 i_4567 (.ZN (n_5207), .A1 (inputB[10]), .A2 (inputA[1]), .A3 (n_5262));
NAND2_X1 i_4566 (.ZN (n_5202), .A1 (n_5212), .A2 (n_5207));
NAND2_X1 i_4565 (.ZN (n_5197), .A1 (inputB[11]), .A2 (inputA[0]));
XOR2_X1 i_4564 (.Z (n_1275), .A (n_5202), .B (n_5197));
OAI21_X1 i_4563 (.ZN (n_5196), .A (n_5261), .B1 (n_5264), .B2 (n_5258));
XOR2_X1 i_4562 (.Z (n_1303), .A (n_1301), .B (n_5196));
AOI21_X1 i_4561 (.ZN (n_5192), .A (n_1257), .B1 (n_1256), .B2 (n_5240));
INV_X1 i_4560 (.ZN (n_1260), .A (n_5192));
AOI21_X1 i_4559 (.ZN (n_5187), .A (n_1252), .B1 (n_1251), .B2 (n_5251));
INV_X1 i_4558 (.ZN (n_5182), .A (n_5187));
XNOR2_X1 i_4556 (.ZN (n_1313), .A (n_1311), .B (n_5187));
AND2_X1 i_4555 (.ZN (n_5181), .A1 (inputB[4]), .A2 (inputA[8]));
NAND2_X1 i_4554 (.ZN (n_5177), .A1 (n_5272), .A2 (n_5181));
AOI22_X1 i_4552 (.ZN (n_5172), .A1 (inputB[3]), .A2 (inputA[8]), .B1 (inputB[4]), .B2 (inputA[7]));
INV_X1 i_4551 (.ZN (n_5171), .A (n_5172));
NAND2_X1 i_4550 (.ZN (n_5167), .A1 (n_5177), .A2 (n_5171));
NAND2_X1 i_4548 (.ZN (n_5163), .A1 (inputB[5]), .A2 (inputA[6]));
XOR2_X1 i_4547 (.Z (n_5162), .A (n_5167), .B (n_5163));
XOR2_X1 i_4546 (.Z (n_1308), .A (n_1306), .B (n_5162));
AOI21_X1 i_4544 (.ZN (n_5161), .A (n_1206), .B1 (n_1205), .B2 (n_5283));
INV_X1 i_4543 (.ZN (n_5160), .A (n_5161));
XNOR2_X1 i_4542 (.ZN (n_5159), .A (n_1261), .B (n_5161));
AOI21_X1 i_4540 (.ZN (n_5158), .A (n_1267), .B1 (n_1266), .B2 (n_5159));
INV_X1 i_4539 (.ZN (n_1270), .A (n_5158));
NAND2_X1 i_4538 (.ZN (n_5156), .A1 (n_5222), .A2 (n_5218));
NAND2_X1 i_4536 (.ZN (n_1283), .A1 (n_5227), .A2 (n_5156));
OAI21_X1 i_4535 (.ZN (n_1276), .A (n_5207), .B1 (n_5217), .B2 (n_5197));
NAND2_X1 i_4534 (.ZN (n_5155), .A1 (inputB[2]), .A2 (inputA[10]));
NAND2_X1 i_4532 (.ZN (n_5154), .A1 (n_5234), .A2 (n_5155));
INV_X1 i_4531 (.ZN (n_5153), .A (n_5154));
OAI21_X1 i_4530 (.ZN (n_5150), .A (n_5154), .B1 (n_5234), .B2 (n_5155));
NAND2_X1 i_4528 (.ZN (n_5149), .A1 (inputB[3]), .A2 (inputA[9]));
XOR2_X1 i_4527 (.Z (n_1351), .A (n_5150), .B (n_5149));
AOI21_X1 i_4526 (.ZN (n_5148), .A (n_5181), .B1 (inputB[5]), .B2 (inputA[7]));
INV_X1 i_4524 (.ZN (n_5147), .A (n_5148));
NAND3_X1 i_4523 (.ZN (n_5146), .A1 (inputB[5]), .A2 (inputA[7]), .A3 (n_5181));
NAND2_X1 i_4522 (.ZN (n_5144), .A1 (n_5147), .A2 (n_5146));
NAND2_X1 i_4520 (.ZN (n_5143), .A1 (inputB[6]), .A2 (inputA[6]));
XOR2_X1 i_4519 (.Z (n_1344), .A (n_5144), .B (n_5143));
AND2_X1 i_4518 (.ZN (n_5142), .A1 (inputB[11]), .A2 (inputA[1]));
AOI21_X1 i_4516 (.ZN (n_5141), .A (n_5142), .B1 (inputB[10]), .B2 (inputA[2]));
INV_X1 i_4515 (.ZN (n_5140), .A (n_5141));
NAND3_X1 i_4514 (.ZN (n_5139), .A1 (inputB[10]), .A2 (inputA[2]), .A3 (n_5142));
NAND2_X1 i_4512 (.ZN (n_5138), .A1 (n_5140), .A2 (n_5139));
NAND2_X1 i_4511 (.ZN (n_5136), .A1 (inputB[12]), .A2 (inputA[0]));
XOR2_X1 i_4510 (.Z (n_1330), .A (n_5138), .B (n_5136));
AOI21_X1 i_4508 (.ZN (n_5135), .A (n_1302), .B1 (n_1301), .B2 (n_5196));
INV_X1 i_4507 (.ZN (n_5134), .A (n_5135));
XNOR2_X1 i_4506 (.ZN (n_1366), .A (n_1364), .B (n_5135));
AOI21_X1 i_4504 (.ZN (n_5133), .A (n_1307), .B1 (n_1306), .B2 (n_5162));
INV_X1 i_4503 (.ZN (n_1310), .A (n_5133));
AOI21_X1 i_4502 (.ZN (n_5132), .A (n_1312), .B1 (n_1311), .B2 (n_5182));
INV_X1 i_4501 (.ZN (n_1315), .A (n_5132));
AOI21_X1 i_4500 (.ZN (n_5129), .A (n_1262), .B1 (n_1261), .B2 (n_5160));
INV_X1 i_4499 (.ZN (n_5128), .A (n_5129));
AOI21_X1 i_4498 (.ZN (n_5127), .A (n_1317), .B1 (n_1316), .B2 (n_5128));
INV_X1 i_4497 (.ZN (n_1320), .A (n_5127));
OAI21_X1 i_4496 (.ZN (n_5126), .A (n_5177), .B1 (n_5172), .B2 (n_5163));
OAI22_X1 i_4495 (.ZN (n_5125), .A1 (n_5279), .A2 (n_5234), .B1 (n_5236), .B2 (n_5232));
NOR2_X1 i_4494 (.ZN (n_5123), .A1 (n_5126), .A2 (n_5125));
NAND2_X1 i_4493 (.ZN (n_5122), .A1 (n_5126), .A2 (n_5125));
OAI21_X1 i_4492 (.ZN (n_5121), .A (n_5122), .B1 (n_5126), .B2 (n_5125));
NAND2_X1 i_4491 (.ZN (n_5120), .A1 (inputB[0]), .A2 (inputA[12]));
XOR2_X1 i_4490 (.Z (n_5119), .A (n_5121), .B (n_5120));
XOR2_X1 i_4489 (.Z (n_1376), .A (n_1374), .B (n_5119));
XNOR2_X1 i_4488 (.ZN (n_5118), .A (n_1316), .B (n_5129));
AOI21_X1 i_4487 (.ZN (n_5117), .A (n_1322), .B1 (n_1321), .B2 (n_5118));
INV_X1 i_4486 (.ZN (n_1325), .A (n_5117));
OAI21_X1 i_4485 (.ZN (n_1345), .A (n_5146), .B1 (n_5148), .B2 (n_5143));
AOI22_X1 i_4484 (.ZN (n_5116), .A1 (inputB[7]), .A2 (inputA[5]), .B1 (inputB[8]), .B2 (inputA[4]));
AND2_X1 i_4483 (.ZN (n_5115), .A1 (inputB[8]), .A2 (inputA[5]));
NAND2_X1 i_4482 (.ZN (n_5113), .A1 (n_5229), .A2 (n_5115));
NAND2_X1 i_4481 (.ZN (n_5111), .A1 (inputB[9]), .A2 (inputA[3]));
OAI21_X1 i_4480 (.ZN (n_1338), .A (n_5113), .B1 (n_5116), .B2 (n_5111));
OAI21_X1 i_4479 (.ZN (n_1359), .A (n_5122), .B1 (n_5123), .B2 (n_5120));
NAND2_X1 i_4478 (.ZN (n_5106), .A1 (inputB[0]), .A2 (inputA[13]));
INV_X1 i_4477 (.ZN (n_5105), .A (n_5106));
AND2_X1 i_4476 (.ZN (n_5102), .A1 (inputB[1]), .A2 (inputA[12]));
XNOR2_X1 i_4475 (.ZN (n_5101), .A (n_5106), .B (n_5102));
OAI22_X1 i_4474 (.ZN (n_5097), .A1 (n_5234), .A2 (n_5155), .B1 (n_5153), .B2 (n_5149));
XOR2_X1 i_4473 (.Z (n_1420), .A (n_5101), .B (n_5097));
AND2_X1 i_4472 (.ZN (n_5096), .A1 (inputB[6]), .A2 (inputA[7]));
AOI21_X1 i_4471 (.ZN (n_5095), .A (n_5096), .B1 (inputB[5]), .B2 (inputA[8]));
INV_X1 i_4470 (.ZN (n_5091), .A (n_5095));
NAND3_X1 i_4469 (.ZN (n_5086), .A1 (inputB[5]), .A2 (inputA[8]), .A3 (n_5096));
NAND2_X1 i_4468 (.ZN (n_5082), .A1 (n_5091), .A2 (n_5086));
NAND2_X1 i_4467 (.ZN (n_5081), .A1 (inputB[7]), .A2 (inputA[6]));
XOR2_X1 i_4466 (.Z (n_1407), .A (n_5082), .B (n_5081));
AOI21_X1 i_4465 (.ZN (n_5076), .A (n_5115), .B1 (inputB[9]), .B2 (inputA[4]));
INV_X1 i_4464 (.ZN (n_5071), .A (n_5076));
NAND3_X1 i_4463 (.ZN (n_5067), .A1 (inputB[9]), .A2 (inputA[4]), .A3 (n_5115));
NAND2_X1 i_4462 (.ZN (n_5066), .A1 (n_5071), .A2 (n_5067));
NAND2_X1 i_4461 (.ZN (n_5061), .A1 (inputB[10]), .A2 (inputA[3]));
XOR2_X1 i_4460 (.Z (n_1400), .A (n_5066), .B (n_5061));
AOI21_X1 i_4459 (.ZN (n_5056), .A (n_1365), .B1 (n_1364), .B2 (n_5134));
INV_X1 i_4458 (.ZN (n_1368), .A (n_5056));
OAI21_X1 i_4457 (.ZN (n_5051), .A (n_5139), .B1 (n_5141), .B2 (n_5136));
XOR2_X1 i_4456 (.Z (n_1429), .A (n_1427), .B (n_5051));
AOI21_X1 i_4455 (.ZN (n_5050), .A (n_1375), .B1 (n_1374), .B2 (n_5119));
INV_X1 i_4454 (.ZN (n_1378), .A (n_5050));
NAND2_X1 i_4453 (.ZN (n_5047), .A1 (inputB[12]), .A2 (inputA[2]));
INV_X1 i_4452 (.ZN (n_5046), .A (n_5047));
NAND2_X1 i_4451 (.ZN (n_5042), .A1 (n_5142), .A2 (n_5046));
AOI22_X1 i_4450 (.ZN (n_5041), .A1 (inputB[11]), .A2 (inputA[2]), .B1 (inputB[12]), .B2 (inputA[1]));
INV_X1 i_4449 (.ZN (n_5040), .A (n_5041));
NAND2_X1 i_4448 (.ZN (n_5038), .A1 (n_5042), .A2 (n_5040));
NAND2_X1 i_4447 (.ZN (n_5037), .A1 (inputB[13]), .A2 (inputA[0]));
XOR2_X1 i_4446 (.Z (n_5036), .A (n_5038), .B (n_5037));
XOR2_X1 i_4445 (.Z (n_1439), .A (n_1437), .B (n_5036));
AOI21_X1 i_4444 (.ZN (n_5035), .A (n_5116), .B1 (n_5229), .B2 (n_5115));
XNOR2_X1 i_4442 (.ZN (n_5034), .A (n_5111), .B (n_5035));
AOI21_X1 i_4441 (.ZN (n_5033), .A (n_1370), .B1 (n_1369), .B2 (n_5034));
INV_X1 i_4440 (.ZN (n_5030), .A (n_5033));
XNOR2_X1 i_4438 (.ZN (n_1444), .A (n_1442), .B (n_5033));
XOR2_X1 i_4437 (.Z (n_5029), .A (n_1369), .B (n_5034));
AOI21_X1 i_4436 (.ZN (n_5028), .A (n_1380), .B1 (n_1379), .B2 (n_5029));
INV_X1 i_4434 (.ZN (n_1383), .A (n_5028));
AND2_X1 i_4433 (.ZN (n_5027), .A1 (inputB[3]), .A2 (inputA[11]));
NAND3_X1 i_4432 (.ZN (n_5026), .A1 (inputB[2]), .A2 (inputA[10]), .A3 (n_5027));
AOI22_X1 i_4430 (.ZN (n_5025), .A1 (inputB[2]), .A2 (inputA[11]), .B1 (inputB[3]), .B2 (inputA[10]));
INV_X1 i_4429 (.ZN (n_5023), .A (n_5025));
NAND2_X1 i_4428 (.ZN (n_5022), .A1 (n_5026), .A2 (n_5023));
NAND2_X1 i_4426 (.ZN (n_5021), .A1 (inputB[4]), .A2 (inputA[9]));
XOR2_X1 i_4425 (.Z (n_5020), .A (n_5022), .B (n_5021));
XOR2_X1 i_4424 (.Z (n_5019), .A (n_1432), .B (n_5020));
XOR2_X1 i_4422 (.Z (n_1449), .A (n_1447), .B (n_5019));
OAI21_X1 i_4421 (.ZN (n_1415), .A (n_5026), .B1 (n_5025), .B2 (n_5021));
OAI21_X1 i_4420 (.ZN (n_1408), .A (n_5086), .B1 (n_5095), .B2 (n_5081));
OAI21_X1 i_4418 (.ZN (n_1394), .A (n_5042), .B1 (n_5041), .B2 (n_5037));
AOI21_X1 i_4417 (.ZN (n_5017), .A (n_1428), .B1 (n_1427), .B2 (n_5051));
INV_X1 i_4416 (.ZN (n_1431), .A (n_5017));
NAND2_X1 i_4414 (.ZN (n_5016), .A1 (inputB[1]), .A2 (inputA[14]));
INV_X1 i_4413 (.ZN (n_5015), .A (n_5016));
NAND2_X1 i_4412 (.ZN (n_5014), .A1 (n_5105), .A2 (n_5015));
AOI22_X1 i_4410 (.ZN (n_5013), .A1 (inputB[1]), .A2 (inputA[13]), .B1 (inputB[0]), .B2 (inputA[14]));
INV_X1 i_4409 (.ZN (n_5012), .A (n_5013));
NAND2_X1 i_4408 (.ZN (n_5009), .A1 (n_5014), .A2 (n_5012));
NAND2_X1 i_4406 (.ZN (n_5008), .A1 (inputB[2]), .A2 (inputA[12]));
XOR2_X1 i_4405 (.Z (n_1489), .A (n_5009), .B (n_5008));
AOI21_X1 i_4404 (.ZN (n_5007), .A (n_5027), .B1 (inputB[4]), .B2 (inputA[10]));
NAND3_X1 i_4402 (.ZN (n_5006), .A1 (inputB[4]), .A2 (inputA[10]), .A3 (n_5027));
INV_X1 i_4401 (.ZN (n_5005), .A (n_5006));
NOR2_X1 i_4400 (.ZN (n_5004), .A1 (n_5007), .A2 (n_5005));
NAND2_X1 i_4398 (.ZN (n_5002), .A1 (inputB[5]), .A2 (inputA[9]));
XNOR2_X1 i_4397 (.ZN (n_1482), .A (n_5004), .B (n_5002));
AOI22_X1 i_4396 (.ZN (n_5001), .A1 (inputB[9]), .A2 (inputA[5]), .B1 (inputB[10]), .B2 (inputA[4]));
INV_X1 i_4394 (.ZN (n_5000), .A (n_5001));
NAND4_X1 i_4393 (.ZN (n_4999), .A1 (inputB[9]), .A2 (inputA[5]), .A3 (inputB[10]), .A4 (inputA[4]));
NAND2_X1 i_4392 (.ZN (n_4998), .A1 (n_5000), .A2 (n_4999));
NAND2_X1 i_4390 (.ZN (n_4997), .A1 (inputB[11]), .A2 (inputA[3]));
XOR2_X1 i_4389 (.Z (n_1468), .A (n_4998), .B (n_4997));
NAND2_X1 i_4388 (.ZN (n_4996), .A1 (inputB[13]), .A2 (inputA[1]));
INV_X1 i_4386 (.ZN (n_4994), .A (n_4996));
NAND2_X1 i_4385 (.ZN (n_4993), .A1 (n_5046), .A2 (n_4994));
NAND2_X1 i_4384 (.ZN (n_4991), .A1 (n_5047), .A2 (n_4996));
AND2_X1 i_4383 (.ZN (n_4986), .A1 (n_4993), .A2 (n_4991));
AND2_X1 i_4382 (.ZN (n_4985), .A1 (inputB[14]), .A2 (inputA[0]));
XOR2_X1 i_4381 (.Z (n_1461), .A (n_4986), .B (n_4985));
AOI21_X1 i_4380 (.ZN (n_4981), .A (n_1438), .B1 (n_1437), .B2 (n_5036));
INV_X1 i_4379 (.ZN (n_1441), .A (n_4981));
AOI21_X1 i_4378 (.ZN (n_4977), .A (n_1433), .B1 (n_1432), .B2 (n_5020));
INV_X1 i_4377 (.ZN (n_1436), .A (n_4977));
AOI21_X1 i_4376 (.ZN (n_4976), .A (n_1443), .B1 (n_1442), .B2 (n_5030));
INV_X1 i_4375 (.ZN (n_1446), .A (n_4976));
OAI21_X1 i_4374 (.ZN (n_4971), .A (n_5067), .B1 (n_5076), .B2 (n_5061));
XOR2_X1 i_4373 (.Z (n_4967), .A (n_1494), .B (n_4971));
XOR2_X1 i_4372 (.Z (n_1511), .A (n_1509), .B (n_4967));
AOI22_X1 i_4371 (.ZN (n_4966), .A1 (n_5105), .A2 (n_5102), .B1 (n_5101), .B2 (n_5097));
INV_X1 i_4370 (.ZN (n_4962), .A (n_4966));
XNOR2_X1 i_4369 (.ZN (n_4961), .A (n_1499), .B (n_4966));
XOR2_X1 i_4368 (.Z (n_1516), .A (n_1514), .B (n_4961));
AOI21_X1 i_4367 (.ZN (n_4957), .A (n_1448), .B1 (n_1447), .B2 (n_5019));
INV_X1 i_4366 (.ZN (n_1451), .A (n_4957));
XOR2_X1 i_4365 (.Z (n_4956), .A (n_1379), .B (n_5029));
AOI21_X1 i_4364 (.ZN (n_4951), .A (n_1385), .B1 (n_1384), .B2 (n_4956));
INV_X1 i_4363 (.ZN (n_4950), .A (n_4951));
AOI21_X1 i_4362 (.ZN (n_4946), .A (n_1453), .B1 (n_1452), .B2 (n_4950));
INV_X1 i_4361 (.ZN (n_1456), .A (n_4946));
AOI22_X1 i_4360 (.ZN (n_4942), .A1 (inputB[6]), .A2 (inputA[8]), .B1 (inputB[7]), .B2 (inputA[7]));
NAND2_X1 i_4359 (.ZN (n_4941), .A1 (inputB[7]), .A2 (inputA[8]));
INV_X1 i_4358 (.ZN (n_4936), .A (n_4941));
NAND2_X1 i_4357 (.ZN (n_4935), .A1 (n_5096), .A2 (n_4936));
NAND2_X1 i_4356 (.ZN (n_4932), .A1 (inputB[8]), .A2 (inputA[6]));
OAI21_X1 i_4355 (.ZN (n_1476), .A (n_4935), .B1 (n_4942), .B2 (n_4932));
OAI21_X1 i_4354 (.ZN (n_1469), .A (n_4999), .B1 (n_5001), .B2 (n_4997));
AOI21_X1 i_4353 (.ZN (n_4931), .A (n_1495), .B1 (n_1494), .B2 (n_4971));
INV_X1 i_4352 (.ZN (n_1498), .A (n_4931));
NAND2_X1 i_4351 (.ZN (n_4926), .A1 (inputB[2]), .A2 (inputA[13]));
INV_X1 i_4350 (.ZN (n_4922), .A (n_4926));
NAND2_X1 i_4349 (.ZN (n_4921), .A1 (n_5015), .A2 (n_4922));
OAI21_X1 i_4348 (.ZN (n_4920), .A (n_4921), .B1 (n_5015), .B2 (n_4922));
NAND2_X1 i_4347 (.ZN (n_4919), .A1 (inputB[3]), .A2 (inputA[12]));
XOR2_X1 i_4346 (.Z (n_1561), .A (n_4920), .B (n_4919));
NAND2_X1 i_4345 (.ZN (n_4916), .A1 (inputB[8]), .A2 (inputA[7]));
INV_X1 i_4344 (.ZN (n_4915), .A (n_4916));
NAND2_X1 i_4343 (.ZN (n_4914), .A1 (n_4936), .A2 (n_4915));
OAI21_X1 i_4342 (.ZN (n_4913), .A (n_4914), .B1 (n_4936), .B2 (n_4915));
NAND2_X1 i_4341 (.ZN (n_4912), .A1 (inputB[9]), .A2 (inputA[6]));
XOR2_X1 i_4340 (.Z (n_1547), .A (n_4913), .B (n_4912));
AND2_X1 i_4339 (.ZN (n_4909), .A1 (inputB[11]), .A2 (inputA[4]));
AOI21_X1 i_4338 (.ZN (n_4908), .A (n_4909), .B1 (inputB[10]), .B2 (inputA[5]));
INV_X1 i_4337 (.ZN (n_4907), .A (n_4908));
NAND3_X1 i_4336 (.ZN (n_4906), .A1 (inputB[10]), .A2 (inputA[5]), .A3 (n_4909));
NAND2_X1 i_4335 (.ZN (n_4905), .A1 (n_4907), .A2 (n_4906));
NAND2_X1 i_4334 (.ZN (n_4904), .A1 (inputB[12]), .A2 (inputA[3]));
XOR2_X1 i_4333 (.Z (n_1540), .A (n_4905), .B (n_4904));
AOI21_X1 i_4332 (.ZN (n_4903), .A (n_1500), .B1 (n_1499), .B2 (n_4962));
INV_X1 i_4331 (.ZN (n_1503), .A (n_4903));
NAND2_X1 i_4330 (.ZN (n_4902), .A1 (n_4991), .A2 (n_4985));
NAND2_X1 i_4329 (.ZN (n_4901), .A1 (n_4993), .A2 (n_4902));
XOR2_X1 i_4328 (.Z (n_1576), .A (n_1574), .B (n_4901));
AOI21_X1 i_4327 (.ZN (n_4900), .A (n_4942), .B1 (n_5096), .B2 (n_4936));
XNOR2_X1 i_4326 (.ZN (n_4899), .A (n_4932), .B (n_4900));
AOI21_X1 i_4324 (.ZN (n_4898), .A (n_1505), .B1 (n_1504), .B2 (n_4899));
INV_X1 i_4323 (.ZN (n_1508), .A (n_4898));
AOI21_X1 i_4322 (.ZN (n_4895), .A (n_1510), .B1 (n_1509), .B2 (n_4967));
INV_X1 i_4320 (.ZN (n_1513), .A (n_4895));
AND2_X1 i_4319 (.ZN (n_4894), .A1 (inputB[5]), .A2 (inputA[10]));
AOI21_X1 i_4318 (.ZN (n_4893), .A (n_4894), .B1 (inputB[4]), .B2 (inputA[11]));
INV_X1 i_4316 (.ZN (n_4892), .A (n_4893));
NAND3_X1 i_4315 (.ZN (n_4891), .A1 (inputB[4]), .A2 (inputA[11]), .A3 (n_4894));
NAND2_X1 i_4314 (.ZN (n_4888), .A1 (n_4892), .A2 (n_4891));
NAND2_X1 i_4312 (.ZN (n_4887), .A1 (inputB[6]), .A2 (inputA[9]));
XOR2_X1 i_4311 (.Z (n_4886), .A (n_4888), .B (n_4887));
XOR2_X1 i_4310 (.Z (n_1581), .A (n_1579), .B (n_4886));
AOI21_X1 i_4308 (.ZN (n_4885), .A (n_1515), .B1 (n_1514), .B2 (n_4961));
INV_X1 i_4307 (.ZN (n_1518), .A (n_4885));
XOR2_X1 i_4306 (.Z (n_4884), .A (n_1504), .B (n_4899));
AOI21_X1 i_4304 (.ZN (n_4883), .A (n_1520), .B1 (n_1519), .B2 (n_4884));
INV_X1 i_4303 (.ZN (n_1523), .A (n_4883));
NAND2_X1 i_4302 (.ZN (n_4882), .A1 (inputB[15]), .A2 (inputA[0]));
AOI22_X1 i_4300 (.ZN (n_4881), .A1 (inputB[13]), .A2 (inputA[2]), .B1 (inputB[14]), .B2 (inputA[1]));
NAND3_X1 i_4299 (.ZN (n_4880), .A1 (inputB[14]), .A2 (inputA[2]), .A3 (n_4994));
INV_X1 i_4298 (.ZN (n_4879), .A (n_4880));
NOR2_X1 i_4296 (.ZN (n_4878), .A1 (n_4881), .A2 (n_4879));
XNOR2_X1 i_4295 (.ZN (n_4877), .A (n_4882), .B (n_4878));
XOR2_X1 i_4294 (.Z (n_4874), .A (n_1584), .B (n_4877));
XOR2_X1 i_4292 (.Z (n_1596), .A (n_1594), .B (n_4874));
XOR2_X1 i_4291 (.Z (n_4873), .A (n_1519), .B (n_4884));
AOI21_X1 i_4290 (.ZN (n_4872), .A (n_1525), .B1 (n_1524), .B2 (n_4873));
INV_X1 i_4288 (.ZN (n_1528), .A (n_4872));
OAI21_X1 i_4287 (.ZN (n_1555), .A (n_4891), .B1 (n_4893), .B2 (n_4887));
AOI22_X1 i_4286 (.ZN (n_1548), .A1 (n_4941), .A2 (n_4916), .B1 (n_4914), .B2 (n_4912));
OAI21_X1 i_4284 (.ZN (n_1534), .A (n_4880), .B1 (n_4882), .B2 (n_4881));
AOI21_X1 i_4283 (.ZN (n_4871), .A (n_1575), .B1 (n_1574), .B2 (n_4901));
INV_X1 i_4282 (.ZN (n_1578), .A (n_4871));
AND2_X1 i_4280 (.ZN (n_4870), .A1 (inputB[0]), .A2 (inputA[16]));
AOI22_X1 i_4279 (.ZN (n_4869), .A1 (n_5016), .A2 (n_4926), .B1 (n_4921), .B2 (n_4919));
NOR2_X1 i_4278 (.ZN (n_4868), .A1 (n_4870), .A2 (n_4869));
NAND2_X1 i_4276 (.ZN (n_4865), .A1 (n_4870), .A2 (n_4869));
OAI21_X1 i_4275 (.ZN (n_4863), .A (n_4865), .B1 (n_4870), .B2 (n_4869));
NAND2_X1 i_4274 (.ZN (n_4858), .A1 (inputB[1]), .A2 (inputA[15]));
XOR2_X1 i_4272 (.Z (n_1647), .A (n_4863), .B (n_4858));
AOI22_X1 i_4271 (.ZN (n_4857), .A1 (inputB[2]), .A2 (inputA[14]), .B1 (inputB[3]), .B2 (inputA[13]));
INV_X1 i_4270 (.ZN (n_4854), .A (n_4857));
AND2_X1 i_4268 (.ZN (n_4853), .A1 (inputB[3]), .A2 (inputA[14]));
NAND2_X1 i_4267 (.ZN (n_4849), .A1 (n_4922), .A2 (n_4853));
NAND2_X1 i_4266 (.ZN (n_4848), .A1 (n_4854), .A2 (n_4849));
NAND2_X1 i_4264 (.ZN (n_4843), .A1 (inputB[4]), .A2 (inputA[12]));
XOR2_X1 i_4263 (.Z (n_1641), .A (n_4848), .B (n_4843));
AOI22_X1 i_4262 (.ZN (n_4842), .A1 (inputB[8]), .A2 (inputA[8]), .B1 (inputB[9]), .B2 (inputA[7]));
INV_X1 i_4261 (.ZN (n_4839), .A (n_4842));
NAND2_X1 i_4260 (.ZN (n_4838), .A1 (inputB[9]), .A2 (inputA[8]));
INV_X1 i_4259 (.ZN (n_4834), .A (n_4838));
NAND2_X1 i_4258 (.ZN (n_4833), .A1 (n_4915), .A2 (n_4834));
NAND2_X1 i_4257 (.ZN (n_4832), .A1 (n_4839), .A2 (n_4833));
NAND2_X1 i_4256 (.ZN (n_4828), .A1 (inputB[10]), .A2 (inputA[6]));
XOR2_X1 i_4255 (.Z (n_1627), .A (n_4832), .B (n_4828));
AOI22_X1 i_4254 (.ZN (n_4823), .A1 (inputB[11]), .A2 (inputA[5]), .B1 (inputB[12]), .B2 (inputA[4]));
INV_X1 i_4253 (.ZN (n_4819), .A (n_4823));
AND2_X1 i_4252 (.ZN (n_4818), .A1 (inputB[12]), .A2 (inputA[5]));
NAND2_X1 i_4251 (.ZN (n_4817), .A1 (n_4909), .A2 (n_4818));
NAND2_X1 i_4250 (.ZN (n_4813), .A1 (n_4819), .A2 (n_4817));
NAND2_X1 i_4249 (.ZN (n_4808), .A1 (inputB[13]), .A2 (inputA[3]));
XOR2_X1 i_4248 (.Z (n_1620), .A (n_4813), .B (n_4808));
OAI21_X1 i_4247 (.ZN (n_4807), .A (n_4906), .B1 (n_4908), .B2 (n_4904));
XOR2_X1 i_4246 (.Z (n_1656), .A (n_1654), .B (n_4807));
AOI21_X1 i_4245 (.ZN (n_4804), .A (n_1585), .B1 (n_1584), .B2 (n_4877));
INV_X1 i_4244 (.ZN (n_1588), .A (n_4804));
AOI21_X1 i_4243 (.ZN (n_4803), .A (n_5013), .B1 (n_5014), .B2 (n_5008));
AOI21_X1 i_4242 (.ZN (n_4802), .A (n_5007), .B1 (n_5006), .B2 (n_5002));
NOR2_X1 i_4241 (.ZN (n_4798), .A1 (n_4803), .A2 (n_4802));
NAND2_X1 i_4240 (.ZN (n_4794), .A1 (n_4803), .A2 (n_4802));
NAND2_X1 i_4239 (.ZN (n_4793), .A1 (inputB[0]), .A2 (inputA[15]));
OAI21_X1 i_4238 (.ZN (n_4789), .A (n_4794), .B1 (n_4798), .B2 (n_4793));
XOR2_X1 i_4237 (.Z (n_1661), .A (n_1659), .B (n_4789));
OAI21_X1 i_4236 (.ZN (n_4788), .A (n_4794), .B1 (n_4803), .B2 (n_4802));
XOR2_X1 i_4235 (.Z (n_4787), .A (n_4793), .B (n_4788));
AOI21_X1 i_4234 (.ZN (n_4786), .A (n_1590), .B1 (n_1589), .B2 (n_4787));
INV_X1 i_4233 (.ZN (n_1593), .A (n_4786));
AND2_X1 i_4232 (.ZN (n_4785), .A1 (inputB[6]), .A2 (inputA[11]));
NAND2_X1 i_4231 (.ZN (n_4784), .A1 (n_4894), .A2 (n_4785));
AOI22_X1 i_4230 (.ZN (n_4783), .A1 (inputB[5]), .A2 (inputA[11]), .B1 (inputB[6]), .B2 (inputA[10]));
INV_X1 i_4229 (.ZN (n_4782), .A (n_4783));
NAND2_X1 i_4228 (.ZN (n_4781), .A1 (n_4784), .A2 (n_4782));
NAND2_X1 i_4227 (.ZN (n_4780), .A1 (inputB[7]), .A2 (inputA[9]));
XOR2_X1 i_4226 (.Z (n_4779), .A (n_4781), .B (n_4780));
XOR2_X1 i_4225 (.Z (n_1666), .A (n_1664), .B (n_4779));
AOI21_X1 i_4224 (.ZN (n_4776), .A (n_1580), .B1 (n_1579), .B2 (n_4886));
INV_X1 i_4223 (.ZN (n_4775), .A (n_4776));
XNOR2_X1 i_4222 (.ZN (n_1676), .A (n_1674), .B (n_4776));
AOI22_X1 i_4221 (.ZN (n_4774), .A1 (inputB[14]), .A2 (inputA[2]), .B1 (inputB[15]), .B2 (inputA[1]));
INV_X1 i_4220 (.ZN (n_4773), .A (n_4774));
AND2_X1 i_4219 (.ZN (n_4772), .A1 (inputB[15]), .A2 (inputA[2]));
NAND3_X1 i_4218 (.ZN (n_4769), .A1 (inputB[14]), .A2 (inputA[1]), .A3 (n_4772));
NAND2_X1 i_4217 (.ZN (n_4768), .A1 (n_4773), .A2 (n_4769));
NAND2_X1 i_4216 (.ZN (n_4767), .A1 (inputB[16]), .A2 (inputA[0]));
XOR2_X1 i_4215 (.Z (n_4766), .A (n_4768), .B (n_4767));
XOR2_X1 i_4214 (.Z (n_4765), .A (n_1669), .B (n_4766));
XOR2_X1 i_4213 (.Z (n_1681), .A (n_1679), .B (n_4765));
XOR2_X1 i_4212 (.Z (n_4764), .A (n_1589), .B (n_4787));
AOI21_X1 i_4211 (.ZN (n_4763), .A (n_1600), .B1 (n_1599), .B2 (n_4764));
INV_X1 i_4210 (.ZN (n_1603), .A (n_4763));
XOR2_X1 i_4209 (.Z (n_4762), .A (n_1599), .B (n_4764));
AOI21_X1 i_4208 (.ZN (n_4761), .A (n_1605), .B1 (n_1604), .B2 (n_4762));
INV_X1 i_4207 (.ZN (n_1608), .A (n_4761));
OAI21_X1 i_4206 (.ZN (n_1642), .A (n_4849), .B1 (n_4857), .B2 (n_4843));
OAI21_X1 i_4205 (.ZN (n_1635), .A (n_4784), .B1 (n_4783), .B2 (n_4780));
OAI21_X1 i_4203 (.ZN (n_1621), .A (n_4817), .B1 (n_4823), .B2 (n_4808));
OAI21_X1 i_4202 (.ZN (n_1614), .A (n_4769), .B1 (n_4774), .B2 (n_4767));
OAI21_X1 i_4201 (.ZN (n_1648), .A (n_4865), .B1 (n_4868), .B2 (n_4858));
AOI22_X1 i_4199 (.ZN (n_4760), .A1 (inputB[0]), .A2 (inputA[17]), .B1 (inputB[1]), .B2 (inputA[16]));
INV_X1 i_4198 (.ZN (n_4759), .A (n_4760));
NAND2_X1 i_4197 (.ZN (n_4758), .A1 (inputB[1]), .A2 (inputA[17]));
INV_X1 i_4195 (.ZN (n_4755), .A (n_4758));
NAND2_X1 i_4194 (.ZN (n_4754), .A1 (n_4870), .A2 (n_4755));
NAND2_X1 i_4193 (.ZN (n_4753), .A1 (n_4759), .A2 (n_4754));
NAND2_X1 i_4191 (.ZN (n_4752), .A1 (inputB[2]), .A2 (inputA[15]));
XOR2_X1 i_4190 (.Z (n_1733), .A (n_4753), .B (n_4752));
AOI21_X1 i_4189 (.ZN (n_4751), .A (n_4785), .B1 (inputB[7]), .B2 (inputA[10]));
INV_X1 i_4187 (.ZN (n_4748), .A (n_4751));
NAND3_X1 i_4186 (.ZN (n_4747), .A1 (inputB[7]), .A2 (inputA[10]), .A3 (n_4785));
NAND2_X1 i_4185 (.ZN (n_4746), .A1 (n_4748), .A2 (n_4747));
NAND2_X1 i_4183 (.ZN (n_4745), .A1 (inputB[8]), .A2 (inputA[9]));
XOR2_X1 i_4182 (.Z (n_1719), .A (n_4746), .B (n_4745));
NAND2_X1 i_4181 (.ZN (n_4744), .A1 (inputB[10]), .A2 (inputA[7]));
INV_X1 i_4179 (.ZN (n_4743), .A (n_4744));
NAND2_X1 i_4178 (.ZN (n_4742), .A1 (n_4834), .A2 (n_4743));
OAI21_X1 i_4177 (.ZN (n_4741), .A (n_4742), .B1 (n_4834), .B2 (n_4743));
NAND2_X1 i_4175 (.ZN (n_4740), .A1 (inputB[11]), .A2 (inputA[6]));
XOR2_X1 i_4174 (.Z (n_1712), .A (n_4741), .B (n_4740));
AOI21_X1 i_4173 (.ZN (n_4739), .A (n_4772), .B1 (inputB[16]), .B2 (inputA[1]));
INV_X1 i_4171 (.ZN (n_4738), .A (n_4739));
NAND3_X1 i_4170 (.ZN (n_4737), .A1 (inputB[16]), .A2 (inputA[1]), .A3 (n_4772));
NAND2_X1 i_4169 (.ZN (n_4736), .A1 (n_4738), .A2 (n_4737));
NAND2_X1 i_4167 (.ZN (n_4735), .A1 (inputB[17]), .A2 (inputA[0]));
XOR2_X1 i_4166 (.Z (n_1698), .A (n_4736), .B (n_4735));
AOI21_X1 i_4165 (.ZN (n_4732), .A (n_1660), .B1 (n_1659), .B2 (n_4789));
INV_X1 i_4163 (.ZN (n_1663), .A (n_4732));
OAI21_X1 i_4162 (.ZN (n_4730), .A (n_4833), .B1 (n_4842), .B2 (n_4828));
XOR2_X1 i_4161 (.Z (n_1740), .A (n_1738), .B (n_4730));
AOI21_X1 i_4159 (.ZN (n_4725), .A (n_1670), .B1 (n_1669), .B2 (n_4766));
INV_X1 i_4158 (.ZN (n_1673), .A (n_4725));
AOI21_X1 i_4157 (.ZN (n_4724), .A (n_1675), .B1 (n_1674), .B2 (n_4775));
INV_X1 i_4155 (.ZN (n_1678), .A (n_4724));
AOI21_X1 i_4154 (.ZN (n_4721), .A (n_4818), .B1 (inputB[13]), .B2 (inputA[4]));
INV_X1 i_4153 (.ZN (n_4720), .A (n_4721));
NAND3_X1 i_4151 (.ZN (n_4715), .A1 (inputB[13]), .A2 (inputA[4]), .A3 (n_4818));
NAND2_X1 i_4150 (.ZN (n_4710), .A1 (n_4720), .A2 (n_4715));
NAND2_X1 i_4149 (.ZN (n_4709), .A1 (inputB[14]), .A2 (inputA[3]));
XOR2_X1 i_4147 (.Z (n_4705), .A (n_4710), .B (n_4709));
XOR2_X1 i_4146 (.Z (n_1755), .A (n_1753), .B (n_4705));
AOI21_X1 i_4145 (.ZN (n_4701), .A (n_1655), .B1 (n_1654), .B2 (n_4807));
INV_X1 i_4143 (.ZN (n_4700), .A (n_4701));
XNOR2_X1 i_4142 (.ZN (n_4699), .A (n_1743), .B (n_4701));
XOR2_X1 i_4141 (.Z (n_1760), .A (n_1758), .B (n_4699));
AOI21_X1 i_4140 (.ZN (n_4695), .A (n_1665), .B1 (n_1664), .B2 (n_4779));
INV_X1 i_4139 (.ZN (n_4694), .A (n_4695));
XNOR2_X1 i_4138 (.ZN (n_1765), .A (n_1763), .B (n_4695));
AOI21_X1 i_4137 (.ZN (n_4690), .A (n_1595), .B1 (n_1594), .B2 (n_4874));
INV_X1 i_4136 (.ZN (n_4685), .A (n_4690));
AOI21_X1 i_4135 (.ZN (n_4681), .A (n_1685), .B1 (n_1684), .B2 (n_4685));
INV_X1 i_4134 (.ZN (n_1688), .A (n_4681));
AOI21_X1 i_4133 (.ZN (n_4680), .A (n_4853), .B1 (inputB[4]), .B2 (inputA[13]));
INV_X1 i_4132 (.ZN (n_4679), .A (n_4680));
NAND3_X1 i_4131 (.ZN (n_4675), .A1 (inputB[4]), .A2 (inputA[13]), .A3 (n_4853));
NAND2_X1 i_4130 (.ZN (n_4670), .A1 (n_4679), .A2 (n_4675));
NAND2_X1 i_4129 (.ZN (n_4666), .A1 (inputB[5]), .A2 (inputA[12]));
XOR2_X1 i_4128 (.Z (n_4665), .A (n_4670), .B (n_4666));
XOR2_X1 i_4127 (.Z (n_4660), .A (n_1748), .B (n_4665));
XOR2_X1 i_4126 (.Z (n_1770), .A (n_1768), .B (n_4660));
XNOR2_X1 i_4125 (.ZN (n_4655), .A (n_1684), .B (n_4690));
AOI21_X1 i_4124 (.ZN (n_4654), .A (n_1690), .B1 (n_1689), .B2 (n_4655));
INV_X1 i_4123 (.ZN (n_1693), .A (n_4654));
OAI21_X1 i_4122 (.ZN (n_1720), .A (n_4747), .B1 (n_4751), .B2 (n_4745));
AOI22_X1 i_4121 (.ZN (n_1713), .A1 (n_4838), .A2 (n_4744), .B1 (n_4742), .B2 (n_4740));
OAI21_X1 i_4120 (.ZN (n_1699), .A (n_4737), .B1 (n_4739), .B2 (n_4735));
AOI21_X1 i_4119 (.ZN (n_4651), .A (n_1739), .B1 (n_1738), .B2 (n_4730));
INV_X1 i_4118 (.ZN (n_1742), .A (n_4651));
AND2_X1 i_4117 (.ZN (n_4650), .A1 (inputB[5]), .A2 (inputA[13]));
AOI21_X1 i_4116 (.ZN (n_4649), .A (n_4650), .B1 (inputB[4]), .B2 (inputA[14]));
INV_X1 i_4115 (.ZN (n_4646), .A (n_4649));
NAND3_X1 i_4114 (.ZN (n_4645), .A1 (inputB[4]), .A2 (inputA[14]), .A3 (n_4650));
NAND2_X1 i_4113 (.ZN (n_4644), .A1 (n_4646), .A2 (n_4645));
NAND2_X1 i_4112 (.ZN (n_4643), .A1 (inputB[6]), .A2 (inputA[12]));
XOR2_X1 i_4111 (.Z (n_1815), .A (n_4644), .B (n_4643));
AOI22_X1 i_4110 (.ZN (n_4642), .A1 (inputB[7]), .A2 (inputA[11]), .B1 (inputB[8]), .B2 (inputA[10]));
INV_X1 i_4109 (.ZN (n_4639), .A (n_4642));
NAND4_X1 i_4108 (.ZN (n_4638), .A1 (inputB[7]), .A2 (inputA[11]), .A3 (inputB[8]), .A4 (inputA[10]));
NAND2_X1 i_4107 (.ZN (n_4637), .A1 (n_4639), .A2 (n_4638));
NAND2_X1 i_4106 (.ZN (n_4636), .A1 (inputB[9]), .A2 (inputA[9]));
XOR2_X1 i_4105 (.Z (n_1808), .A (n_4637), .B (n_4636));
AND2_X1 i_4104 (.ZN (n_4635), .A1 (inputB[14]), .A2 (inputA[4]));
AOI21_X1 i_4103 (.ZN (n_4634), .A (n_4635), .B1 (inputB[13]), .B2 (inputA[5]));
INV_X1 i_4102 (.ZN (n_4633), .A (n_4634));
NAND3_X1 i_4101 (.ZN (n_4632), .A1 (inputB[13]), .A2 (inputA[5]), .A3 (n_4635));
NAND2_X1 i_4100 (.ZN (n_4631), .A1 (n_4633), .A2 (n_4632));
NAND2_X1 i_4099 (.ZN (n_4630), .A1 (inputB[15]), .A2 (inputA[3]));
XOR2_X1 i_4098 (.Z (n_1794), .A (n_4631), .B (n_4630));
AOI22_X1 i_4097 (.ZN (n_4629), .A1 (inputB[16]), .A2 (inputA[2]), .B1 (inputB[17]), .B2 (inputA[1]));
INV_X1 i_4096 (.ZN (n_4628), .A (n_4629));
NAND4_X1 i_4095 (.ZN (n_4625), .A1 (inputB[16]), .A2 (inputA[2]), .A3 (inputB[17]), .A4 (inputA[1]));
NAND2_X1 i_4094 (.ZN (n_4624), .A1 (n_4628), .A2 (n_4625));
NAND2_X1 i_4093 (.ZN (n_4623), .A1 (inputB[18]), .A2 (inputA[0]));
XOR2_X1 i_4092 (.Z (n_1787), .A (n_4624), .B (n_4623));
OAI21_X1 i_4091 (.ZN (n_4622), .A (n_4715), .B1 (n_4721), .B2 (n_4709));
XOR2_X1 i_4090 (.Z (n_1837), .A (n_1835), .B (n_4622));
OAI21_X1 i_4089 (.ZN (n_4621), .A (n_4754), .B1 (n_4760), .B2 (n_4752));
OAI21_X1 i_4088 (.ZN (n_4618), .A (n_4675), .B1 (n_4680), .B2 (n_4666));
OR2_X1 i_4087 (.ZN (n_4617), .A1 (n_4621), .A2 (n_4618));
NAND2_X1 i_4086 (.ZN (n_4616), .A1 (n_4621), .A2 (n_4618));
AND2_X1 i_4085 (.ZN (n_4615), .A1 (n_4617), .A2 (n_4616));
AND2_X1 i_4084 (.ZN (n_4614), .A1 (inputB[0]), .A2 (inputA[18]));
XOR2_X1 i_4083 (.Z (n_1829), .A (n_4615), .B (n_4614));
AOI21_X1 i_4082 (.ZN (n_4613), .A (n_1749), .B1 (n_1748), .B2 (n_4665));
INV_X1 i_4081 (.ZN (n_1752), .A (n_4613));
NAND2_X1 i_4080 (.ZN (n_4612), .A1 (inputB[2]), .A2 (inputA[16]));
INV_X1 i_4079 (.ZN (n_4611), .A (n_4612));
NAND2_X1 i_4078 (.ZN (n_4610), .A1 (n_4755), .A2 (n_4611));
OAI21_X1 i_4077 (.ZN (n_4609), .A (n_4610), .B1 (n_4755), .B2 (n_4611));
NAND2_X1 i_4076 (.ZN (n_4608), .A1 (inputB[3]), .A2 (inputA[15]));
XOR2_X1 i_4074 (.Z (n_4607), .A (n_4609), .B (n_4608));
XOR2_X1 i_4073 (.Z (n_1842), .A (n_1840), .B (n_4607));
AOI21_X1 i_4072 (.ZN (n_4604), .A (n_1759), .B1 (n_1758), .B2 (n_4699));
INV_X1 i_4070 (.ZN (n_1762), .A (n_4604));
AOI21_X1 i_4069 (.ZN (n_4603), .A (n_1744), .B1 (n_1743), .B2 (n_4700));
INV_X1 i_4068 (.ZN (n_4602), .A (n_4603));
XNOR2_X1 i_4066 (.ZN (n_1852), .A (n_1850), .B (n_4603));
AOI21_X1 i_4065 (.ZN (n_4601), .A (n_1754), .B1 (n_1753), .B2 (n_4705));
INV_X1 i_4064 (.ZN (n_4600), .A (n_4601));
XNOR2_X1 i_4062 (.ZN (n_1857), .A (n_1855), .B (n_4601));
AOI21_X1 i_4061 (.ZN (n_4599), .A (n_1769), .B1 (n_1768), .B2 (n_4660));
INV_X1 i_4060 (.ZN (n_1772), .A (n_4599));
AOI21_X1 i_4058 (.ZN (n_4598), .A (n_1680), .B1 (n_1679), .B2 (n_4765));
INV_X1 i_4057 (.ZN (n_4595), .A (n_4598));
AOI21_X1 i_4056 (.ZN (n_4593), .A (n_1774), .B1 (n_1773), .B2 (n_4595));
INV_X1 i_4054 (.ZN (n_1777), .A (n_4593));
AOI22_X1 i_4053 (.ZN (n_4588), .A1 (inputB[10]), .A2 (inputA[8]), .B1 (inputB[11]), .B2 (inputA[7]));
NAND3_X1 i_4052 (.ZN (n_4587), .A1 (inputB[11]), .A2 (inputA[8]), .A3 (n_4743));
INV_X1 i_4050 (.ZN (n_4584), .A (n_4587));
NOR2_X1 i_4049 (.ZN (n_4583), .A1 (n_4588), .A2 (n_4584));
NAND2_X1 i_4048 (.ZN (n_4578), .A1 (inputB[12]), .A2 (inputA[6]));
XNOR2_X1 i_4046 (.ZN (n_4573), .A (n_4583), .B (n_4578));
XOR2_X1 i_4045 (.Z (n_4568), .A (n_1845), .B (n_4573));
XOR2_X1 i_4044 (.Z (n_1867), .A (n_1865), .B (n_4568));
XNOR2_X1 i_4042 (.ZN (n_4563), .A (n_1773), .B (n_4598));
AOI21_X1 i_4041 (.ZN (n_4562), .A (n_1779), .B1 (n_1778), .B2 (n_4563));
INV_X1 i_4040 (.ZN (n_1782), .A (n_4562));
AOI21_X1 i_4038 (.ZN (n_4559), .A (n_1764), .B1 (n_1763), .B2 (n_4694));
INV_X1 i_4037 (.ZN (n_4558), .A (n_4559));
XNOR2_X1 i_4036 (.ZN (n_4553), .A (n_1860), .B (n_4559));
XOR2_X1 i_4034 (.Z (n_4552), .A (n_1870), .B (n_4553));
XOR2_X1 i_4033 (.Z (n_1877), .A (n_1875), .B (n_4552));
OAI21_X1 i_4032 (.ZN (n_1816), .A (n_4645), .B1 (n_4649), .B2 (n_4643));
OAI21_X1 i_4030 (.ZN (n_1809), .A (n_4638), .B1 (n_4642), .B2 (n_4636));
OAI21_X1 i_4029 (.ZN (n_1795), .A (n_4632), .B1 (n_4634), .B2 (n_4630));
OAI21_X1 i_4028 (.ZN (n_1788), .A (n_4625), .B1 (n_4629), .B2 (n_4623));
NAND2_X1 i_4026 (.ZN (n_4548), .A1 (n_4617), .A2 (n_4614));
NAND2_X1 i_4025 (.ZN (n_1830), .A1 (n_4616), .A2 (n_4548));
AND2_X1 i_4024 (.ZN (n_4543), .A1 (inputB[1]), .A2 (inputA[19]));
AOI22_X1 i_4022 (.ZN (n_4538), .A1 (inputB[1]), .A2 (inputA[18]), .B1 (inputB[0]), .B2 (inputA[19]));
AOI21_X1 i_4021 (.ZN (n_4537), .A (n_4538), .B1 (n_4614), .B2 (n_4543));
AOI22_X1 i_4020 (.ZN (n_4534), .A1 (n_4758), .A2 (n_4612), .B1 (n_4610), .B2 (n_4608));
XOR2_X1 i_4018 (.Z (n_1925), .A (n_4537), .B (n_4534));
AOI22_X1 i_4017 (.ZN (n_4533), .A1 (inputB[5]), .A2 (inputA[14]), .B1 (inputB[6]), .B2 (inputA[13]));
INV_X1 i_4016 (.ZN (n_4529), .A (n_4533));
NAND3_X1 i_4014 (.ZN (n_4528), .A1 (inputB[6]), .A2 (inputA[14]), .A3 (n_4650));
NAND2_X1 i_4013 (.ZN (n_4523), .A1 (n_4529), .A2 (n_4528));
NAND2_X1 i_4012 (.ZN (n_4518), .A1 (inputB[7]), .A2 (inputA[12]));
XOR2_X1 i_4010 (.Z (n_1912), .A (n_4523), .B (n_4518));
AND2_X1 i_4009 (.ZN (n_4517), .A1 (inputB[9]), .A2 (inputA[10]));
AOI21_X1 i_4008 (.ZN (n_4514), .A (n_4517), .B1 (inputB[8]), .B2 (inputA[11]));
INV_X1 i_4007 (.ZN (n_4513), .A (n_4514));
NAND3_X1 i_4006 (.ZN (n_4512), .A1 (inputB[8]), .A2 (inputA[11]), .A3 (n_4517));
NAND2_X1 i_4005 (.ZN (n_4511), .A1 (n_4513), .A2 (n_4512));
NAND2_X1 i_4004 (.ZN (n_4510), .A1 (inputB[10]), .A2 (inputA[9]));
XOR2_X1 i_4003 (.Z (n_1905), .A (n_4511), .B (n_4510));
AOI22_X1 i_4002 (.ZN (n_4509), .A1 (inputB[14]), .A2 (inputA[5]), .B1 (inputB[15]), .B2 (inputA[4]));
INV_X1 i_4001 (.ZN (n_4508), .A (n_4509));
NAND3_X1 i_4000 (.ZN (n_4507), .A1 (inputB[15]), .A2 (inputA[5]), .A3 (n_4635));
NAND2_X1 i_3999 (.ZN (n_4506), .A1 (n_4508), .A2 (n_4507));
NAND2_X1 i_3998 (.ZN (n_4505), .A1 (inputB[16]), .A2 (inputA[3]));
XOR2_X1 i_3997 (.Z (n_1891), .A (n_4506), .B (n_4505));
AND2_X1 i_3996 (.ZN (n_4504), .A1 (inputB[18]), .A2 (inputA[1]));
AOI21_X1 i_3995 (.ZN (n_4501), .A (n_4504), .B1 (inputB[17]), .B2 (inputA[2]));
INV_X1 i_3994 (.ZN (n_4500), .A (n_4501));
NAND3_X1 i_3993 (.ZN (n_4499), .A1 (inputB[17]), .A2 (inputA[2]), .A3 (n_4504));
NAND2_X1 i_3992 (.ZN (n_4498), .A1 (n_4500), .A2 (n_4499));
NAND2_X1 i_3991 (.ZN (n_4497), .A1 (inputB[19]), .A2 (inputA[0]));
XOR2_X1 i_3990 (.Z (n_1884), .A (n_4498), .B (n_4497));
AOI21_X1 i_3989 (.ZN (n_4496), .A (n_4588), .B1 (n_4587), .B2 (n_4578));
XOR2_X1 i_3988 (.Z (n_1934), .A (n_1932), .B (n_4496));
AOI21_X1 i_3987 (.ZN (n_4494), .A (n_1846), .B1 (n_1845), .B2 (n_4573));
INV_X1 i_3986 (.ZN (n_1849), .A (n_4494));
AOI21_X1 i_3985 (.ZN (n_4493), .A (n_1851), .B1 (n_1850), .B2 (n_4602));
INV_X1 i_3984 (.ZN (n_1854), .A (n_4493));
AOI21_X1 i_3983 (.ZN (n_4492), .A (n_1856), .B1 (n_1855), .B2 (n_4600));
INV_X1 i_3982 (.ZN (n_1859), .A (n_4492));
NAND2_X1 i_3981 (.ZN (n_4491), .A1 (inputB[13]), .A2 (inputA[6]));
AOI22_X1 i_3980 (.ZN (n_4490), .A1 (inputB[11]), .A2 (inputA[8]), .B1 (inputB[12]), .B2 (inputA[7]));
NAND2_X1 i_3979 (.ZN (n_4488), .A1 (inputB[12]), .A2 (inputA[8]));
INV_X1 i_3978 (.ZN (n_4487), .A (n_4488));
NAND3_X1 i_3977 (.ZN (n_4486), .A1 (inputB[11]), .A2 (inputA[7]), .A3 (n_4487));
INV_X1 i_3976 (.ZN (n_4485), .A (n_4486));
NOR2_X1 i_3975 (.ZN (n_4484), .A1 (n_4490), .A2 (n_4485));
XNOR2_X1 i_3974 (.ZN (n_4483), .A (n_4491), .B (n_4484));
XOR2_X1 i_3973 (.Z (n_1949), .A (n_1947), .B (n_4483));
NAND2_X1 i_3972 (.ZN (n_4480), .A1 (inputB[3]), .A2 (inputA[17]));
INV_X1 i_3971 (.ZN (n_4479), .A (n_4480));
NAND2_X1 i_3970 (.ZN (n_4478), .A1 (n_4611), .A2 (n_4479));
AOI22_X1 i_3969 (.ZN (n_4477), .A1 (inputB[2]), .A2 (inputA[17]), .B1 (inputB[3]), .B2 (inputA[16]));
INV_X1 i_3968 (.ZN (n_4476), .A (n_4477));
NAND2_X1 i_3967 (.ZN (n_4475), .A1 (n_4478), .A2 (n_4476));
NAND2_X1 i_3966 (.ZN (n_4473), .A1 (inputB[4]), .A2 (inputA[15]));
XOR2_X1 i_3965 (.Z (n_4472), .A (n_4475), .B (n_4473));
XOR2_X1 i_3964 (.Z (n_1944), .A (n_1942), .B (n_4472));
AOI21_X1 i_3963 (.ZN (n_4471), .A (n_1841), .B1 (n_1840), .B2 (n_4607));
INV_X1 i_3962 (.ZN (n_4470), .A (n_4471));
XNOR2_X1 i_3961 (.ZN (n_1959), .A (n_1957), .B (n_4471));
AOI21_X1 i_3960 (.ZN (n_4469), .A (n_1866), .B1 (n_1865), .B2 (n_4568));
INV_X1 i_3959 (.ZN (n_1869), .A (n_4469));
AOI21_X1 i_3958 (.ZN (n_4467), .A (n_1861), .B1 (n_1860), .B2 (n_4558));
INV_X1 i_3957 (.ZN (n_4466), .A (n_4467));
XNOR2_X1 i_3956 (.ZN (n_1969), .A (n_1967), .B (n_4467));
AOI21_X1 i_3955 (.ZN (n_4465), .A (n_1871), .B1 (n_1870), .B2 (n_4553));
INV_X1 i_3954 (.ZN (n_1874), .A (n_4465));
AOI21_X1 i_3953 (.ZN (n_4464), .A (n_1876), .B1 (n_1875), .B2 (n_4552));
INV_X1 i_3952 (.ZN (n_1879), .A (n_4464));
AOI21_X1 i_3951 (.ZN (n_4463), .A (n_1836), .B1 (n_1835), .B2 (n_4622));
INV_X1 i_3950 (.ZN (n_4462), .A (n_4463));
XNOR2_X1 i_3949 (.ZN (n_4459), .A (n_1937), .B (n_4463));
XOR2_X1 i_3948 (.Z (n_4458), .A (n_1952), .B (n_4459));
XOR2_X1 i_3947 (.Z (n_4457), .A (n_1962), .B (n_4458));
XOR2_X1 i_3946 (.Z (n_4456), .A (n_1972), .B (n_4457));
XOR2_X1 i_3945 (.Z (n_1979), .A (n_1977), .B (n_4456));
OAI21_X1 i_3944 (.ZN (n_1920), .A (n_4478), .B1 (n_4477), .B2 (n_4473));
OAI21_X1 i_3943 (.ZN (n_1913), .A (n_4528), .B1 (n_4533), .B2 (n_4518));
OAI21_X1 i_3941 (.ZN (n_1899), .A (n_4486), .B1 (n_4491), .B2 (n_4490));
OAI21_X1 i_3940 (.ZN (n_1892), .A (n_4507), .B1 (n_4509), .B2 (n_4505));
AOI21_X1 i_3939 (.ZN (n_4455), .A (n_1933), .B1 (n_1932), .B2 (n_4496));
INV_X1 i_3937 (.ZN (n_1936), .A (n_4455));
AOI22_X1 i_3936 (.ZN (n_4454), .A1 (n_4614), .A2 (n_4543), .B1 (n_4537), .B2 (n_4534));
INV_X1 i_3935 (.ZN (n_1926), .A (n_4454));
NAND2_X1 i_3933 (.ZN (n_4453), .A1 (inputB[4]), .A2 (inputA[16]));
INV_X1 i_3932 (.ZN (n_4452), .A (n_4453));
NAND2_X1 i_3931 (.ZN (n_4450), .A1 (n_4480), .A2 (n_4453));
AOI22_X1 i_3929 (.ZN (n_4448), .A1 (n_4479), .A2 (n_4452), .B1 (n_4480), .B2 (n_4453));
AND2_X1 i_3928 (.ZN (n_4443), .A1 (inputB[5]), .A2 (inputA[15]));
XOR2_X1 i_3927 (.Z (n_2021), .A (n_4448), .B (n_4443));
AOI22_X1 i_3925 (.ZN (n_4442), .A1 (inputB[6]), .A2 (inputA[14]), .B1 (inputB[7]), .B2 (inputA[13]));
INV_X1 i_3924 (.ZN (n_4439), .A (n_4442));
NAND2_X1 i_3923 (.ZN (n_4438), .A1 (inputB[7]), .A2 (inputA[14]));
INV_X1 i_3921 (.ZN (n_4434), .A (n_4438));
NAND3_X1 i_3920 (.ZN (n_4433), .A1 (inputB[6]), .A2 (inputA[13]), .A3 (n_4434));
NAND2_X1 i_3919 (.ZN (n_4428), .A1 (n_4439), .A2 (n_4433));
NAND2_X1 i_3917 (.ZN (n_4423), .A1 (inputB[8]), .A2 (inputA[12]));
XOR2_X1 i_3916 (.Z (n_2014), .A (n_4428), .B (n_4423));
NAND2_X1 i_3915 (.ZN (n_4418), .A1 (inputB[13]), .A2 (inputA[7]));
INV_X1 i_3913 (.ZN (n_4417), .A (n_4418));
NAND2_X1 i_3912 (.ZN (n_4413), .A1 (n_4487), .A2 (n_4417));
NAND2_X1 i_3911 (.ZN (n_4408), .A1 (n_4488), .A2 (n_4418));
AND2_X1 i_3909 (.ZN (n_4404), .A1 (n_4413), .A2 (n_4408));
AND2_X1 i_3908 (.ZN (n_4403), .A1 (inputB[14]), .A2 (inputA[6]));
XOR2_X1 i_3907 (.Z (n_2000), .A (n_4404), .B (n_4403));
AOI22_X1 i_3905 (.ZN (n_4398), .A1 (inputB[15]), .A2 (inputA[5]), .B1 (inputB[16]), .B2 (inputA[4]));
INV_X1 i_3904 (.ZN (n_4397), .A (n_4398));
NAND4_X1 i_3903 (.ZN (n_4393), .A1 (inputB[15]), .A2 (inputA[4]), .A3 (inputB[16]), .A4 (inputA[5]));
NAND2_X1 i_3901 (.ZN (n_4389), .A1 (n_4397), .A2 (n_4393));
NAND2_X1 i_3900 (.ZN (n_4388), .A1 (inputB[17]), .A2 (inputA[3]));
XOR2_X1 i_3899 (.Z (n_1993), .A (n_4389), .B (n_4388));
AOI21_X1 i_3897 (.ZN (n_4384), .A (n_1938), .B1 (n_1937), .B2 (n_4462));
INV_X1 i_3896 (.ZN (n_1941), .A (n_4384));
OAI21_X1 i_3895 (.ZN (n_4383), .A (n_4499), .B1 (n_4501), .B2 (n_4497));
XOR2_X1 i_3893 (.Z (n_2040), .A (n_2038), .B (n_4383));
AOI21_X1 i_3892 (.ZN (n_4382), .A (n_1948), .B1 (n_1947), .B2 (n_4483));
INV_X1 i_3891 (.ZN (n_1951), .A (n_4382));
AOI21_X1 i_3889 (.ZN (n_4379), .A (n_1943), .B1 (n_1942), .B2 (n_4472));
INV_X1 i_3888 (.ZN (n_1946), .A (n_4379));
AOI21_X1 i_3887 (.ZN (n_4378), .A (n_1958), .B1 (n_1957), .B2 (n_4470));
INV_X1 i_3885 (.ZN (n_1961), .A (n_4378));
AOI21_X1 i_3884 (.ZN (n_4373), .A (n_1953), .B1 (n_1952), .B2 (n_4459));
INV_X1 i_3883 (.ZN (n_1956), .A (n_4373));
AND2_X1 i_3881 (.ZN (n_4372), .A1 (inputB[10]), .A2 (inputA[11]));
NAND2_X1 i_3880 (.ZN (n_4368), .A1 (n_4517), .A2 (n_4372));
AOI22_X1 i_3879 (.ZN (n_4364), .A1 (inputB[9]), .A2 (inputA[11]), .B1 (inputB[10]), .B2 (inputA[10]));
INV_X1 i_3877 (.ZN (n_4363), .A (n_4364));
NAND2_X1 i_3876 (.ZN (n_4362), .A1 (n_4368), .A2 (n_4363));
NAND2_X1 i_3875 (.ZN (n_4361), .A1 (inputB[11]), .A2 (inputA[9]));
XOR2_X1 i_3873 (.Z (n_4360), .A (n_4362), .B (n_4361));
XOR2_X1 i_3872 (.Z (n_2050), .A (n_2048), .B (n_4360));
AOI21_X1 i_3871 (.ZN (n_4359), .A (n_4543), .B1 (inputB[0]), .B2 (inputA[20]));
INV_X1 i_3870 (.ZN (n_4357), .A (n_4359));
NAND3_X1 i_3869 (.ZN (n_4356), .A1 (inputB[0]), .A2 (inputA[20]), .A3 (n_4543));
NAND2_X1 i_3868 (.ZN (n_4355), .A1 (n_4357), .A2 (n_4356));
NAND2_X1 i_3867 (.ZN (n_4354), .A1 (inputB[2]), .A2 (inputA[18]));
XOR2_X1 i_3866 (.Z (n_4351), .A (n_4355), .B (n_4354));
XOR2_X1 i_3865 (.Z (n_4350), .A (n_2043), .B (n_4351));
XOR2_X1 i_3864 (.Z (n_2065), .A (n_2063), .B (n_4350));
AOI21_X1 i_3863 (.ZN (n_4349), .A (n_1963), .B1 (n_1962), .B2 (n_4458));
INV_X1 i_3862 (.ZN (n_1966), .A (n_4349));
AOI21_X1 i_3861 (.ZN (n_4348), .A (n_1968), .B1 (n_1967), .B2 (n_4466));
INV_X1 i_3860 (.ZN (n_1971), .A (n_4348));
AOI21_X1 i_3859 (.ZN (n_4347), .A (n_1973), .B1 (n_1972), .B2 (n_4457));
INV_X1 i_3858 (.ZN (n_1976), .A (n_4347));
OAI21_X1 i_3857 (.ZN (n_4345), .A (n_4512), .B1 (n_4514), .B2 (n_4510));
XOR2_X1 i_3856 (.Z (n_4344), .A (n_2033), .B (n_4345));
XOR2_X1 i_3855 (.Z (n_4343), .A (n_2058), .B (n_4344));
XOR2_X1 i_3854 (.Z (n_2075), .A (n_2073), .B (n_4343));
AOI21_X1 i_3853 (.ZN (n_4342), .A (n_1978), .B1 (n_1977), .B2 (n_4456));
INV_X1 i_3852 (.ZN (n_1981), .A (n_4342));
OAI21_X1 i_3851 (.ZN (n_2015), .A (n_4433), .B1 (n_4442), .B2 (n_4423));
OAI21_X1 i_3850 (.ZN (n_2008), .A (n_4368), .B1 (n_4364), .B2 (n_4361));
OAI21_X1 i_3849 (.ZN (n_1994), .A (n_4393), .B1 (n_4398), .B2 (n_4388));
AOI22_X1 i_3848 (.ZN (n_4341), .A1 (inputB[18]), .A2 (inputA[2]), .B1 (inputB[19]), .B2 (inputA[1]));
AND2_X1 i_3847 (.ZN (n_4340), .A1 (inputB[19]), .A2 (inputA[2]));
NAND2_X1 i_3846 (.ZN (n_4339), .A1 (n_4504), .A2 (n_4340));
NAND2_X1 i_3845 (.ZN (n_4337), .A1 (inputB[20]), .A2 (inputA[0]));
OAI21_X1 i_3844 (.ZN (n_1987), .A (n_4339), .B1 (n_4341), .B2 (n_4337));
AOI21_X1 i_3843 (.ZN (n_4336), .A (n_2034), .B1 (n_2033), .B2 (n_4345));
INV_X1 i_3842 (.ZN (n_2037), .A (n_4336));
NAND2_X1 i_3841 (.ZN (n_4335), .A1 (inputB[2]), .A2 (inputA[20]));
INV_X1 i_3840 (.ZN (n_4334), .A (n_4335));
NAND2_X1 i_3839 (.ZN (n_4333), .A1 (n_4543), .A2 (n_4334));
AOI22_X1 i_3838 (.ZN (n_4330), .A1 (inputB[1]), .A2 (inputA[20]), .B1 (inputB[2]), .B2 (inputA[19]));
INV_X1 i_3837 (.ZN (n_4329), .A (n_4330));
NAND2_X1 i_3836 (.ZN (n_4328), .A1 (n_4333), .A2 (n_4329));
NAND2_X1 i_3835 (.ZN (n_4327), .A1 (inputB[3]), .A2 (inputA[18]));
XOR2_X1 i_3834 (.Z (n_2134), .A (n_4328), .B (n_4327));
NAND2_X1 i_3833 (.ZN (n_4326), .A1 (inputB[8]), .A2 (inputA[13]));
INV_X1 i_3832 (.ZN (n_4324), .A (n_4326));
NAND2_X1 i_3831 (.ZN (n_4323), .A1 (n_4434), .A2 (n_4324));
OAI21_X1 i_3830 (.ZN (n_4322), .A (n_4323), .B1 (n_4434), .B2 (n_4324));
NAND2_X1 i_3829 (.ZN (n_4321), .A1 (inputB[9]), .A2 (inputA[12]));
XOR2_X1 i_3828 (.Z (n_2120), .A (n_4322), .B (n_4321));
AOI21_X1 i_3827 (.ZN (n_4320), .A (n_4372), .B1 (inputB[11]), .B2 (inputA[10]));
INV_X1 i_3826 (.ZN (n_4319), .A (n_4320));
NAND3_X1 i_3825 (.ZN (n_4318), .A1 (inputB[11]), .A2 (inputA[10]), .A3 (n_4372));
NAND2_X1 i_3824 (.ZN (n_4316), .A1 (n_4319), .A2 (n_4318));
NAND2_X1 i_3823 (.ZN (n_4315), .A1 (inputB[12]), .A2 (inputA[9]));
XOR2_X1 i_3822 (.Z (n_2113), .A (n_4316), .B (n_4315));
AOI22_X1 i_3821 (.ZN (n_4314), .A1 (inputB[16]), .A2 (inputA[5]), .B1 (inputB[17]), .B2 (inputA[4]));
INV_X1 i_3820 (.ZN (n_4313), .A (n_4314));
AND2_X1 i_3819 (.ZN (n_4312), .A1 (inputB[17]), .A2 (inputA[5]));
NAND3_X1 i_3818 (.ZN (n_4309), .A1 (inputB[16]), .A2 (inputA[4]), .A3 (n_4312));
NAND2_X1 i_3817 (.ZN (n_4308), .A1 (n_4313), .A2 (n_4309));
NAND2_X1 i_3816 (.ZN (n_4307), .A1 (inputB[18]), .A2 (inputA[3]));
XOR2_X1 i_3815 (.Z (n_2099), .A (n_4308), .B (n_4307));
AOI21_X1 i_3814 (.ZN (n_4306), .A (n_4340), .B1 (inputB[20]), .B2 (inputA[1]));
INV_X1 i_3813 (.ZN (n_4305), .A (n_4306));
NAND3_X1 i_3812 (.ZN (n_4304), .A1 (inputB[20]), .A2 (inputA[1]), .A3 (n_4340));
NAND2_X1 i_3811 (.ZN (n_4303), .A1 (n_4305), .A2 (n_4304));
NAND2_X1 i_3810 (.ZN (n_4301), .A1 (inputB[21]), .A2 (inputA[0]));
XOR2_X1 i_3809 (.Z (n_2092), .A (n_4303), .B (n_4301));
NAND2_X1 i_3808 (.ZN (n_4300), .A1 (n_4408), .A2 (n_4403));
NAND2_X1 i_3807 (.ZN (n_4298), .A1 (n_4413), .A2 (n_4300));
XOR2_X1 i_3805 (.Z (n_2149), .A (n_2147), .B (n_4298));
OAI21_X1 i_3804 (.ZN (n_4293), .A (n_4356), .B1 (n_4359), .B2 (n_4354));
INV_X1 i_3803 (.ZN (n_4292), .A (n_4293));
AOI22_X1 i_3801 (.ZN (n_4289), .A1 (n_4479), .A2 (n_4452), .B1 (n_4450), .B2 (n_4443));
NOR2_X1 i_3800 (.ZN (n_4288), .A1 (n_4292), .A2 (n_4289));
AOI21_X1 i_3799 (.ZN (n_4284), .A (n_4288), .B1 (n_4292), .B2 (n_4289));
AND2_X1 i_3797 (.ZN (n_4283), .A1 (inputB[0]), .A2 (inputA[21]));
XOR2_X1 i_3796 (.Z (n_2141), .A (n_4284), .B (n_4283));
AOI21_X1 i_3795 (.ZN (n_4282), .A (n_2049), .B1 (n_2048), .B2 (n_4360));
INV_X1 i_3793 (.ZN (n_2052), .A (n_4282));
AOI21_X1 i_3792 (.ZN (n_4278), .A (n_2044), .B1 (n_2043), .B2 (n_4351));
INV_X1 i_3791 (.ZN (n_2047), .A (n_4278));
AOI21_X1 i_3789 (.ZN (n_4273), .A (n_2039), .B1 (n_2038), .B2 (n_4383));
INV_X1 i_3788 (.ZN (n_4269), .A (n_4273));
XNOR2_X1 i_3787 (.ZN (n_4268), .A (n_2152), .B (n_4273));
XOR2_X1 i_3785 (.Z (n_2169), .A (n_2167), .B (n_4268));
AND2_X1 i_3784 (.ZN (n_4264), .A1 (inputB[14]), .A2 (inputA[8]));
NAND2_X1 i_3783 (.ZN (n_4263), .A1 (n_4417), .A2 (n_4264));
AOI22_X1 i_3781 (.ZN (n_4262), .A1 (inputB[13]), .A2 (inputA[8]), .B1 (inputB[14]), .B2 (inputA[7]));
INV_X1 i_3780 (.ZN (n_4258), .A (n_4262));
NAND2_X1 i_3779 (.ZN (n_4253), .A1 (n_4263), .A2 (n_4258));
NAND2_X1 i_3777 (.ZN (n_4248), .A1 (inputB[15]), .A2 (inputA[6]));
XOR2_X1 i_3776 (.Z (n_4247), .A (n_4253), .B (n_4248));
XOR2_X1 i_3775 (.Z (n_2164), .A (n_2162), .B (n_4247));
AOI21_X1 i_3773 (.ZN (n_4243), .A (n_2064), .B1 (n_2063), .B2 (n_4350));
INV_X1 i_3772 (.ZN (n_2067), .A (n_4243));
AOI21_X1 i_3771 (.ZN (n_4239), .A (n_2059), .B1 (n_2058), .B2 (n_4344));
INV_X1 i_3769 (.ZN (n_4238), .A (n_4239));
XNOR2_X1 i_3768 (.ZN (n_2179), .A (n_2177), .B (n_4239));
AOI21_X1 i_3767 (.ZN (n_4233), .A (n_4341), .B1 (n_4504), .B2 (n_4340));
XNOR2_X1 i_3765 (.ZN (n_4228), .A (n_4337), .B (n_4233));
XOR2_X1 i_3764 (.Z (n_4223), .A (n_2053), .B (n_4228));
AOI21_X1 i_3763 (.ZN (n_4218), .A (n_2069), .B1 (n_2068), .B2 (n_4223));
INV_X1 i_3761 (.ZN (n_2072), .A (n_4218));
AOI21_X1 i_3760 (.ZN (n_4214), .A (n_2074), .B1 (n_2073), .B2 (n_4343));
INV_X1 i_3759 (.ZN (n_2077), .A (n_4214));
XOR2_X1 i_3757 (.Z (n_4213), .A (n_2068), .B (n_4223));
AOI21_X1 i_3756 (.ZN (n_4212), .A (n_2079), .B1 (n_2078), .B2 (n_4213));
INV_X1 i_3755 (.ZN (n_2082), .A (n_4212));
AOI21_X1 i_3753 (.ZN (n_4209), .A (n_2054), .B1 (n_2053), .B2 (n_4228));
INV_X1 i_3752 (.ZN (n_4208), .A (n_4209));
XNOR2_X1 i_3751 (.ZN (n_4207), .A (n_2172), .B (n_4209));
XOR2_X1 i_3749 (.Z (n_2189), .A (n_2187), .B (n_4207));
XOR2_X1 i_3748 (.Z (n_4205), .A (n_2078), .B (n_4213));
AOI21_X1 i_3747 (.ZN (n_4204), .A (n_2084), .B1 (n_2083), .B2 (n_4205));
INV_X1 i_3745 (.ZN (n_2087), .A (n_4204));
NAND2_X1 i_3744 (.ZN (n_4203), .A1 (inputB[5]), .A2 (inputA[17]));
INV_X1 i_3743 (.ZN (n_4202), .A (n_4203));
NAND2_X1 i_3741 (.ZN (n_4201), .A1 (n_4452), .A2 (n_4202));
AOI22_X1 i_3740 (.ZN (n_4200), .A1 (inputB[4]), .A2 (inputA[17]), .B1 (inputB[5]), .B2 (inputA[16]));
INV_X1 i_3739 (.ZN (n_4197), .A (n_4200));
NAND2_X1 i_3737 (.ZN (n_4196), .A1 (n_4201), .A2 (n_4197));
NAND2_X1 i_3736 (.ZN (n_4195), .A1 (inputB[6]), .A2 (inputA[15]));
XOR2_X1 i_3735 (.Z (n_4194), .A (n_4196), .B (n_4195));
XOR2_X1 i_3734 (.Z (n_4193), .A (n_2157), .B (n_4194));
XOR2_X1 i_3733 (.Z (n_4192), .A (n_2182), .B (n_4193));
XOR2_X1 i_3732 (.Z (n_4190), .A (n_2192), .B (n_4192));
XOR2_X1 i_3731 (.Z (n_2199), .A (n_2197), .B (n_4190));
OAI21_X1 i_3730 (.ZN (n_2128), .A (n_4201), .B1 (n_4200), .B2 (n_4195));
AOI22_X1 i_3729 (.ZN (n_2121), .A1 (n_4438), .A2 (n_4326), .B1 (n_4323), .B2 (n_4321));
OAI21_X1 i_3728 (.ZN (n_2107), .A (n_4263), .B1 (n_4262), .B2 (n_4248));
OAI21_X1 i_3727 (.ZN (n_2100), .A (n_4309), .B1 (n_4314), .B2 (n_4307));
AOI21_X1 i_3726 (.ZN (n_4189), .A (n_2148), .B1 (n_2147), .B2 (n_4298));
INV_X1 i_3725 (.ZN (n_2151), .A (n_4189));
NOR2_X1 i_3724 (.ZN (n_4188), .A1 (n_4288), .A2 (n_4283));
AOI21_X1 i_3723 (.ZN (n_2142), .A (n_4188), .B1 (n_4292), .B2 (n_4289));
NAND2_X1 i_3722 (.ZN (n_4187), .A1 (inputB[3]), .A2 (inputA[19]));
INV_X1 i_3721 (.ZN (n_4186), .A (n_4187));
NAND2_X1 i_3720 (.ZN (n_4184), .A1 (n_4334), .A2 (n_4186));
NAND2_X1 i_3719 (.ZN (n_4183), .A1 (n_4335), .A2 (n_4187));
AND2_X1 i_3718 (.ZN (n_4182), .A1 (n_4184), .A2 (n_4183));
AND2_X1 i_3717 (.ZN (n_4181), .A1 (inputB[4]), .A2 (inputA[18]));
XOR2_X1 i_3716 (.Z (n_2248), .A (n_4182), .B (n_4181));
NAND2_X1 i_3715 (.ZN (n_4180), .A1 (inputB[6]), .A2 (inputA[16]));
INV_X1 i_3714 (.ZN (n_4179), .A (n_4180));
NAND2_X1 i_3713 (.ZN (n_4176), .A1 (n_4202), .A2 (n_4179));
OAI21_X1 i_3712 (.ZN (n_4175), .A (n_4176), .B1 (n_4202), .B2 (n_4179));
NAND2_X1 i_3711 (.ZN (n_4174), .A1 (inputB[7]), .A2 (inputA[15]));
XOR2_X1 i_3710 (.Z (n_2241), .A (n_4175), .B (n_4174));
AND2_X1 i_3709 (.ZN (n_4173), .A1 (inputB[12]), .A2 (inputA[10]));
AOI21_X1 i_3708 (.ZN (n_4172), .A (n_4173), .B1 (inputB[11]), .B2 (inputA[11]));
INV_X1 i_3707 (.ZN (n_4171), .A (n_4172));
NAND3_X1 i_3706 (.ZN (n_4169), .A1 (inputB[11]), .A2 (inputA[11]), .A3 (n_4173));
NAND2_X1 i_3705 (.ZN (n_4168), .A1 (n_4171), .A2 (n_4169));
NAND2_X1 i_3704 (.ZN (n_4167), .A1 (inputB[13]), .A2 (inputA[9]));
XOR2_X1 i_3703 (.Z (n_2227), .A (n_4168), .B (n_4167));
AOI21_X1 i_3702 (.ZN (n_4166), .A (n_4264), .B1 (inputB[15]), .B2 (inputA[7]));
INV_X1 i_3701 (.ZN (n_4165), .A (n_4166));
NAND3_X1 i_3700 (.ZN (n_4163), .A1 (inputB[15]), .A2 (inputA[7]), .A3 (n_4264));
NAND2_X1 i_3699 (.ZN (n_4162), .A1 (n_4165), .A2 (n_4163));
NAND2_X1 i_3698 (.ZN (n_4161), .A1 (inputB[16]), .A2 (inputA[6]));
XOR2_X1 i_3697 (.Z (n_2220), .A (n_4162), .B (n_4161));
AOI22_X1 i_3696 (.ZN (n_4160), .A1 (inputB[20]), .A2 (inputA[2]), .B1 (inputB[21]), .B2 (inputA[1]));
INV_X1 i_3695 (.ZN (n_4159), .A (n_4160));
NAND4_X1 i_3694 (.ZN (n_4158), .A1 (inputB[20]), .A2 (inputA[2]), .A3 (inputB[21]), .A4 (inputA[1]));
NAND2_X1 i_3693 (.ZN (n_4155), .A1 (n_4159), .A2 (n_4158));
NAND2_X1 i_3692 (.ZN (n_4154), .A1 (inputB[22]), .A2 (inputA[0]));
XOR2_X1 i_3691 (.Z (n_2206), .A (n_4155), .B (n_4154));
AOI21_X1 i_3690 (.ZN (n_4153), .A (n_2153), .B1 (n_2152), .B2 (n_4269));
INV_X1 i_3689 (.ZN (n_2156), .A (n_4153));
OAI21_X1 i_3688 (.ZN (n_4152), .A (n_4318), .B1 (n_4320), .B2 (n_4315));
XOR2_X1 i_3687 (.Z (n_2263), .A (n_2261), .B (n_4152));
AOI21_X1 i_3686 (.ZN (n_4151), .A (n_2163), .B1 (n_2162), .B2 (n_4247));
INV_X1 i_3685 (.ZN (n_2166), .A (n_4151));
AOI21_X1 i_3684 (.ZN (n_4150), .A (n_4330), .B1 (n_4333), .B2 (n_4327));
INV_X1 i_3683 (.ZN (n_4149), .A (n_4150));
AOI22_X1 i_3682 (.ZN (n_4148), .A1 (inputB[0]), .A2 (inputA[22]), .B1 (inputB[1]), .B2 (inputA[21]));
AND2_X1 i_3681 (.ZN (n_4146), .A1 (inputB[1]), .A2 (inputA[22]));
NAND2_X1 i_3680 (.ZN (n_4144), .A1 (n_4283), .A2 (n_4146));
AOI21_X1 i_3679 (.ZN (n_2255), .A (n_4148), .B1 (n_4149), .B2 (n_4144));
OAI21_X1 i_3678 (.ZN (n_4139), .A (n_2255), .B1 (n_4149), .B2 (n_4144));
INV_X1 i_3677 (.ZN (n_4138), .A (n_4139));
AOI21_X1 i_3676 (.ZN (n_4134), .A (n_4138), .B1 (n_4149), .B2 (n_4148));
XOR2_X1 i_3675 (.Z (n_2273), .A (n_2271), .B (n_4134));
AOI21_X1 i_3674 (.ZN (n_4130), .A (n_2173), .B1 (n_2172), .B2 (n_4208));
INV_X1 i_3673 (.ZN (n_2176), .A (n_4130));
AOI21_X1 i_3672 (.ZN (n_4129), .A (n_4312), .B1 (inputB[18]), .B2 (inputA[4]));
INV_X1 i_3671 (.ZN (n_4124), .A (n_4129));
NAND3_X1 i_3670 (.ZN (n_4119), .A1 (inputB[18]), .A2 (inputA[4]), .A3 (n_4312));
NAND2_X1 i_3669 (.ZN (n_4115), .A1 (n_4124), .A2 (n_4119));
NAND2_X1 i_3668 (.ZN (n_4114), .A1 (inputB[19]), .A2 (inputA[3]));
XOR2_X1 i_3667 (.Z (n_4110), .A (n_4115), .B (n_4114));
XOR2_X1 i_3666 (.Z (n_2283), .A (n_2281), .B (n_4110));
NAND2_X1 i_3665 (.ZN (n_4109), .A1 (inputB[9]), .A2 (inputA[14]));
INV_X1 i_3664 (.ZN (n_4105), .A (n_4109));
NAND2_X1 i_3663 (.ZN (n_4104), .A1 (n_4324), .A2 (n_4105));
AOI22_X1 i_3661 (.ZN (n_4099), .A1 (inputB[8]), .A2 (inputA[14]), .B1 (inputB[9]), .B2 (inputA[13]));
INV_X1 i_3660 (.ZN (n_4094), .A (n_4099));
NAND2_X1 i_3659 (.ZN (n_4089), .A1 (n_4104), .A2 (n_4094));
NAND2_X1 i_3657 (.ZN (n_4084), .A1 (inputB[10]), .A2 (inputA[12]));
XOR2_X1 i_3656 (.Z (n_4080), .A (n_4089), .B (n_4084));
XOR2_X1 i_3655 (.Z (n_2278), .A (n_2276), .B (n_4080));
AOI21_X1 i_3653 (.ZN (n_4079), .A (n_2178), .B1 (n_2177), .B2 (n_4238));
INV_X1 i_3652 (.ZN (n_2181), .A (n_4079));
AOI21_X1 i_3651 (.ZN (n_4078), .A (n_2158), .B1 (n_2157), .B2 (n_4194));
INV_X1 i_3649 (.ZN (n_4075), .A (n_4078));
XNOR2_X1 i_3648 (.ZN (n_2293), .A (n_2291), .B (n_4078));
AOI21_X1 i_3647 (.ZN (n_4074), .A (n_2168), .B1 (n_2167), .B2 (n_4268));
INV_X1 i_3645 (.ZN (n_4069), .A (n_4074));
XNOR2_X1 i_3644 (.ZN (n_2298), .A (n_2296), .B (n_4074));
AOI21_X1 i_3643 (.ZN (n_4068), .A (n_2188), .B1 (n_2187), .B2 (n_4207));
INV_X1 i_3641 (.ZN (n_2191), .A (n_4068));
AOI21_X1 i_3640 (.ZN (n_4065), .A (n_2183), .B1 (n_2182), .B2 (n_4193));
INV_X1 i_3639 (.ZN (n_4064), .A (n_4065));
XNOR2_X1 i_3637 (.ZN (n_2308), .A (n_2306), .B (n_4065));
AOI21_X1 i_3636 (.ZN (n_4059), .A (n_2193), .B1 (n_2192), .B2 (n_4192));
INV_X1 i_3635 (.ZN (n_2196), .A (n_4059));
AOI21_X1 i_3633 (.ZN (n_4055), .A (n_2198), .B1 (n_2197), .B2 (n_4190));
INV_X1 i_3632 (.ZN (n_2201), .A (n_4055));
OAI21_X1 i_3631 (.ZN (n_4054), .A (n_4304), .B1 (n_4306), .B2 (n_4301));
XOR2_X1 i_3629 (.Z (n_4053), .A (n_2266), .B (n_4054));
XOR2_X1 i_3628 (.Z (n_4052), .A (n_2286), .B (n_4053));
XOR2_X1 i_3627 (.Z (n_4049), .A (n_2301), .B (n_4052));
XOR2_X1 i_3625 (.Z (n_4048), .A (n_2311), .B (n_4049));
XOR2_X1 i_3624 (.Z (n_2318), .A (n_2316), .B (n_4048));
NAND2_X1 i_3623 (.ZN (n_4047), .A1 (n_4183), .A2 (n_4181));
NAND2_X1 i_3621 (.ZN (n_2249), .A1 (n_4184), .A2 (n_4047));
AOI22_X1 i_3620 (.ZN (n_2242), .A1 (n_4203), .A2 (n_4180), .B1 (n_4176), .B2 (n_4174));
OAI21_X1 i_3619 (.ZN (n_2228), .A (n_4169), .B1 (n_4172), .B2 (n_4167));
OAI21_X1 i_3617 (.ZN (n_2221), .A (n_4163), .B1 (n_4166), .B2 (n_4161));
OAI21_X1 i_3616 (.ZN (n_2207), .A (n_4158), .B1 (n_4160), .B2 (n_4154));
AOI21_X1 i_3615 (.ZN (n_4046), .A (n_2267), .B1 (n_2266), .B2 (n_4054));
INV_X1 i_3613 (.ZN (n_2270), .A (n_4046));
AND3_X1 i_3612 (.ZN (n_4045), .A1 (inputB[0]), .A2 (inputA[23]), .A3 (n_4146));
AOI21_X1 i_3611 (.ZN (n_4042), .A (n_4146), .B1 (inputB[0]), .B2 (inputA[23]));
INV_X1 i_3609 (.ZN (n_4041), .A (n_4042));
NOR2_X1 i_3608 (.ZN (n_4040), .A1 (n_4045), .A2 (n_4042));
AND2_X1 i_3607 (.ZN (n_4039), .A1 (inputB[2]), .A2 (inputA[21]));
XOR2_X1 i_3605 (.Z (n_2374), .A (n_4040), .B (n_4039));
AOI22_X1 i_3604 (.ZN (n_4038), .A1 (inputB[6]), .A2 (inputA[17]), .B1 (inputB[7]), .B2 (inputA[16]));
INV_X1 i_3603 (.ZN (n_4037), .A (n_4038));
NAND3_X1 i_3601 (.ZN (n_4036), .A1 (inputB[7]), .A2 (inputA[17]), .A3 (n_4179));
NAND2_X1 i_3600 (.ZN (n_4035), .A1 (n_4037), .A2 (n_4036));
NAND2_X1 i_3599 (.ZN (n_4034), .A1 (inputB[8]), .A2 (inputA[15]));
XOR2_X1 i_3597 (.Z (n_2360), .A (n_4035), .B (n_4034));
NAND2_X1 i_3596 (.ZN (n_4033), .A1 (inputB[10]), .A2 (inputA[13]));
INV_X1 i_3595 (.ZN (n_4032), .A (n_4033));
NAND2_X1 i_3593 (.ZN (n_4031), .A1 (n_4105), .A2 (n_4032));
NAND2_X1 i_3592 (.ZN (n_4028), .A1 (n_4109), .A2 (n_4033));
AND2_X1 i_3591 (.ZN (n_4027), .A1 (n_4031), .A2 (n_4028));
AND2_X1 i_3589 (.ZN (n_4026), .A1 (inputB[11]), .A2 (inputA[12]));
XOR2_X1 i_3588 (.Z (n_2353), .A (n_4027), .B (n_4026));
AOI22_X1 i_3587 (.ZN (n_4025), .A1 (inputB[15]), .A2 (inputA[8]), .B1 (inputB[16]), .B2 (inputA[7]));
INV_X1 i_3586 (.ZN (n_4024), .A (n_4025));
NAND4_X1 i_3585 (.ZN (n_4021), .A1 (inputB[15]), .A2 (inputA[8]), .A3 (inputB[16]), .A4 (inputA[7]));
NAND2_X1 i_3584 (.ZN (n_4020), .A1 (n_4024), .A2 (n_4021));
NAND2_X1 i_3583 (.ZN (n_4019), .A1 (inputB[17]), .A2 (inputA[6]));
XOR2_X1 i_3582 (.Z (n_2339), .A (n_4020), .B (n_4019));
AND2_X1 i_3581 (.ZN (n_4018), .A1 (inputB[19]), .A2 (inputA[4]));
AOI21_X1 i_3580 (.ZN (n_4017), .A (n_4018), .B1 (inputB[18]), .B2 (inputA[5]));
INV_X1 i_3579 (.ZN (n_4016), .A (n_4017));
NAND3_X1 i_3578 (.ZN (n_4015), .A1 (inputB[18]), .A2 (inputA[5]), .A3 (n_4018));
NAND2_X1 i_3577 (.ZN (n_4014), .A1 (n_4016), .A2 (n_4015));
NAND2_X1 i_3576 (.ZN (n_4013), .A1 (inputB[20]), .A2 (inputA[3]));
XOR2_X1 i_3575 (.Z (n_2332), .A (n_4014), .B (n_4013));
OAI21_X1 i_3574 (.ZN (n_4012), .A (n_4119), .B1 (n_4129), .B2 (n_4114));
XOR2_X1 i_3573 (.Z (n_2386), .A (n_2384), .B (n_4012));
AOI21_X1 i_3572 (.ZN (n_4011), .A (n_4099), .B1 (n_4104), .B2 (n_4084));
XOR2_X1 i_3571 (.Z (n_2381), .A (n_2379), .B (n_4011));
AOI21_X1 i_3570 (.ZN (n_4010), .A (n_2277), .B1 (n_2276), .B2 (n_4080));
INV_X1 i_3569 (.ZN (n_2280), .A (n_4010));
AOI21_X1 i_3568 (.ZN (n_4007), .A (n_2272), .B1 (n_2271), .B2 (n_4134));
INV_X1 i_3567 (.ZN (n_2275), .A (n_4007));
AOI21_X1 i_3566 (.ZN (n_4006), .A (n_2292), .B1 (n_2291), .B2 (n_4075));
INV_X1 i_3565 (.ZN (n_2295), .A (n_4006));
AOI21_X1 i_3564 (.ZN (n_4005), .A (n_2287), .B1 (n_2286), .B2 (n_4053));
INV_X1 i_3563 (.ZN (n_2290), .A (n_4005));
AND2_X1 i_3562 (.ZN (n_4004), .A1 (inputB[13]), .A2 (inputA[11]));
NAND2_X1 i_3561 (.ZN (n_4003), .A1 (n_4173), .A2 (n_4004));
AOI22_X1 i_3560 (.ZN (n_4000), .A1 (inputB[12]), .A2 (inputA[11]), .B1 (inputB[13]), .B2 (inputA[10]));
INV_X1 i_3559 (.ZN (n_3999), .A (n_4000));
NAND2_X1 i_3558 (.ZN (n_3998), .A1 (n_4003), .A2 (n_3999));
NAND2_X1 i_3557 (.ZN (n_3997), .A1 (inputB[14]), .A2 (inputA[9]));
XOR2_X1 i_3556 (.Z (n_3996), .A (n_3998), .B (n_3997));
XOR2_X1 i_3555 (.Z (n_2401), .A (n_2399), .B (n_3996));
NAND2_X1 i_3554 (.ZN (n_3995), .A1 (inputB[4]), .A2 (inputA[20]));
INV_X1 i_3553 (.ZN (n_3994), .A (n_3995));
NAND2_X1 i_3552 (.ZN (n_3993), .A1 (n_4186), .A2 (n_3994));
AOI22_X1 i_3551 (.ZN (n_3992), .A1 (inputB[3]), .A2 (inputA[20]), .B1 (inputB[4]), .B2 (inputA[19]));
INV_X1 i_3550 (.ZN (n_3991), .A (n_3992));
NAND2_X1 i_3549 (.ZN (n_3990), .A1 (n_3993), .A2 (n_3991));
NAND2_X1 i_3548 (.ZN (n_3989), .A1 (inputB[5]), .A2 (inputA[18]));
XOR2_X1 i_3547 (.Z (n_3988), .A (n_3990), .B (n_3989));
XOR2_X1 i_3546 (.Z (n_2396), .A (n_2394), .B (n_3988));
AOI21_X1 i_3545 (.ZN (n_3987), .A (n_2262), .B1 (n_2261), .B2 (n_4152));
INV_X1 i_3544 (.ZN (n_3984), .A (n_3987));
XNOR2_X1 i_3543 (.ZN (n_3982), .A (n_2389), .B (n_3987));
XOR2_X1 i_3542 (.Z (n_2416), .A (n_2414), .B (n_3982));
AOI21_X1 i_3541 (.ZN (n_3977), .A (n_2282), .B1 (n_2281), .B2 (n_4110));
INV_X1 i_3540 (.ZN (n_3976), .A (n_3977));
XNOR2_X1 i_3539 (.ZN (n_2411), .A (n_2409), .B (n_3977));
AOI22_X1 i_3538 (.ZN (n_3973), .A1 (inputB[21]), .A2 (inputA[2]), .B1 (inputB[22]), .B2 (inputA[1]));
INV_X1 i_3537 (.ZN (n_3972), .A (n_3973));
NAND4_X1 i_3536 (.ZN (n_3968), .A1 (inputB[21]), .A2 (inputA[2]), .A3 (inputB[22]), .A4 (inputA[1]));
NAND2_X1 i_3535 (.ZN (n_3967), .A1 (n_3972), .A2 (n_3968));
NAND2_X1 i_3534 (.ZN (n_3962), .A1 (inputB[23]), .A2 (inputA[0]));
XOR2_X1 i_3533 (.Z (n_3958), .A (n_3967), .B (n_3962));
XOR2_X1 i_3532 (.Z (n_3957), .A (n_2404), .B (n_3958));
XOR2_X1 i_3531 (.Z (n_2421), .A (n_2419), .B (n_3957));
AOI21_X1 i_3530 (.ZN (n_3956), .A (n_2307), .B1 (n_2306), .B2 (n_4064));
INV_X1 i_3529 (.ZN (n_2310), .A (n_3956));
AOI21_X1 i_3528 (.ZN (n_3953), .A (n_2302), .B1 (n_2301), .B2 (n_4052));
INV_X1 i_3527 (.ZN (n_3952), .A (n_3953));
XNOR2_X1 i_3526 (.ZN (n_2431), .A (n_2429), .B (n_3953));
AOI21_X1 i_3525 (.ZN (n_3947), .A (n_2312), .B1 (n_2311), .B2 (n_4049));
INV_X1 i_3524 (.ZN (n_2315), .A (n_3947));
AOI21_X1 i_3523 (.ZN (n_3943), .A (n_2317), .B1 (n_2316), .B2 (n_4048));
INV_X1 i_3522 (.ZN (n_2320), .A (n_3943));
AOI21_X1 i_3521 (.ZN (n_3942), .A (n_2297), .B1 (n_2296), .B2 (n_4069));
INV_X1 i_3520 (.ZN (n_3937), .A (n_3942));
XNOR2_X1 i_3519 (.ZN (n_3936), .A (n_2424), .B (n_3942));
XOR2_X1 i_3518 (.Z (n_3933), .A (n_2434), .B (n_3936));
XOR2_X1 i_3517 (.Z (n_2441), .A (n_2439), .B (n_3933));
OAI21_X1 i_3516 (.ZN (n_2361), .A (n_4036), .B1 (n_4038), .B2 (n_4034));
NAND2_X1 i_3515 (.ZN (n_3932), .A1 (n_4028), .A2 (n_4026));
NAND2_X1 i_3513 (.ZN (n_2354), .A1 (n_4031), .A2 (n_3932));
OAI21_X1 i_3512 (.ZN (n_2340), .A (n_4021), .B1 (n_4025), .B2 (n_4019));
OAI21_X1 i_3511 (.ZN (n_2333), .A (n_4015), .B1 (n_4017), .B2 (n_4013));
AOI21_X1 i_3509 (.ZN (n_3928), .A (n_2385), .B1 (n_2384), .B2 (n_4012));
INV_X1 i_3508 (.ZN (n_2388), .A (n_3928));
AOI21_X1 i_3507 (.ZN (n_3927), .A (n_2380), .B1 (n_2379), .B2 (n_4011));
INV_X1 i_3505 (.ZN (n_2383), .A (n_3927));
NAND2_X1 i_3504 (.ZN (n_3922), .A1 (inputB[5]), .A2 (inputA[19]));
INV_X1 i_3503 (.ZN (n_3917), .A (n_3922));
NAND2_X1 i_3501 (.ZN (n_3916), .A1 (n_3994), .A2 (n_3917));
OAI21_X1 i_3500 (.ZN (n_3913), .A (n_3916), .B1 (n_3994), .B2 (n_3917));
NAND2_X1 i_3499 (.ZN (n_3912), .A1 (inputB[6]), .A2 (inputA[18]));
XOR2_X1 i_3497 (.Z (n_2490), .A (n_3913), .B (n_3912));
AOI22_X1 i_3496 (.ZN (n_3911), .A1 (inputB[7]), .A2 (inputA[17]), .B1 (inputB[8]), .B2 (inputA[16]));
INV_X1 i_3495 (.ZN (n_3907), .A (n_3911));
NAND2_X1 i_3493 (.ZN (n_3902), .A1 (inputB[8]), .A2 (inputA[17]));
INV_X1 i_3492 (.ZN (n_3897), .A (n_3902));
NAND3_X1 i_3491 (.ZN (n_3896), .A1 (inputB[7]), .A2 (inputA[16]), .A3 (n_3897));
NAND2_X1 i_3489 (.ZN (n_3893), .A1 (n_3907), .A2 (n_3896));
NAND2_X1 i_3488 (.ZN (n_3892), .A1 (inputB[9]), .A2 (inputA[15]));
XOR2_X1 i_3487 (.Z (n_2483), .A (n_3893), .B (n_3892));
AOI21_X1 i_3485 (.ZN (n_3888), .A (n_4004), .B1 (inputB[14]), .B2 (inputA[10]));
INV_X1 i_3484 (.ZN (n_3887), .A (n_3888));
NAND3_X1 i_3483 (.ZN (n_3886), .A1 (inputB[14]), .A2 (inputA[10]), .A3 (n_4004));
NAND2_X1 i_3481 (.ZN (n_3885), .A1 (n_3887), .A2 (n_3886));
NAND2_X1 i_3480 (.ZN (n_3884), .A1 (inputB[15]), .A2 (inputA[9]));
XOR2_X1 i_3479 (.Z (n_2469), .A (n_3885), .B (n_3884));
AOI22_X1 i_3477 (.ZN (n_3883), .A1 (inputB[16]), .A2 (inputA[8]), .B1 (inputB[17]), .B2 (inputA[7]));
INV_X1 i_3476 (.ZN (n_3882), .A (n_3883));
NAND4_X1 i_3475 (.ZN (n_3881), .A1 (inputB[16]), .A2 (inputA[8]), .A3 (inputB[17]), .A4 (inputA[7]));
NAND2_X1 i_3473 (.ZN (n_3880), .A1 (n_3882), .A2 (n_3881));
NAND2_X1 i_3472 (.ZN (n_3879), .A1 (inputB[18]), .A2 (inputA[6]));
XOR2_X1 i_3471 (.Z (n_2462), .A (n_3880), .B (n_3879));
AOI22_X1 i_3469 (.ZN (n_3878), .A1 (inputB[22]), .A2 (inputA[2]), .B1 (inputB[23]), .B2 (inputA[1]));
INV_X1 i_3468 (.ZN (n_3875), .A (n_3878));
NAND4_X1 i_3467 (.ZN (n_3874), .A1 (inputB[22]), .A2 (inputA[2]), .A3 (inputB[23]), .A4 (inputA[1]));
NAND2_X1 i_3465 (.ZN (n_3873), .A1 (n_3875), .A2 (n_3874));
NAND2_X1 i_3464 (.ZN (n_3872), .A1 (inputB[24]), .A2 (inputA[0]));
XOR2_X1 i_3463 (.Z (n_2448), .A (n_3873), .B (n_3872));
AOI21_X1 i_3461 (.ZN (n_3871), .A (n_2390), .B1 (n_2389), .B2 (n_3984));
INV_X1 i_3460 (.ZN (n_2393), .A (n_3871));
OAI21_X1 i_3459 (.ZN (n_3868), .A (n_4003), .B1 (n_4000), .B2 (n_3997));
XOR2_X1 i_3457 (.Z (n_2512), .A (n_2510), .B (n_3868));
OAI21_X1 i_3456 (.ZN (n_3867), .A (n_3993), .B1 (n_3992), .B2 (n_3989));
INV_X1 i_3455 (.ZN (n_3866), .A (n_3867));
AOI21_X1 i_3453 (.ZN (n_3865), .A (n_4045), .B1 (n_4041), .B2 (n_4039));
NOR2_X1 i_3452 (.ZN (n_3864), .A1 (n_3866), .A2 (n_3865));
AOI21_X1 i_3451 (.ZN (n_3863), .A (n_3864), .B1 (n_3866), .B2 (n_3865));
AND2_X1 i_3449 (.ZN (n_3862), .A1 (inputB[0]), .A2 (inputA[24]));
XOR2_X1 i_3448 (.Z (n_2504), .A (n_3863), .B (n_3862));
AOI21_X1 i_3447 (.ZN (n_3861), .A (n_2400), .B1 (n_2399), .B2 (n_3996));
INV_X1 i_3445 (.ZN (n_2403), .A (n_3861));
AOI21_X1 i_3444 (.ZN (n_3860), .A (n_2395), .B1 (n_2394), .B2 (n_3988));
INV_X1 i_3443 (.ZN (n_2398), .A (n_3860));
AOI21_X1 i_3441 (.ZN (n_3859), .A (n_2410), .B1 (n_2409), .B2 (n_3976));
INV_X1 i_3440 (.ZN (n_2413), .A (n_3859));
AOI22_X1 i_3439 (.ZN (n_3858), .A1 (inputB[19]), .A2 (inputA[5]), .B1 (inputB[20]), .B2 (inputA[4]));
INV_X1 i_3438 (.ZN (n_3857), .A (n_3858));
NAND3_X1 i_3437 (.ZN (n_3854), .A1 (inputB[20]), .A2 (inputA[5]), .A3 (n_4018));
NAND2_X1 i_3436 (.ZN (n_3853), .A1 (n_3857), .A2 (n_3854));
NAND2_X1 i_3435 (.ZN (n_3852), .A1 (inputB[21]), .A2 (inputA[3]));
XOR2_X1 i_3434 (.Z (n_3851), .A (n_3853), .B (n_3852));
XOR2_X1 i_3433 (.Z (n_2532), .A (n_2530), .B (n_3851));
OAI21_X1 i_3432 (.ZN (n_3850), .A (n_3968), .B1 (n_3973), .B2 (n_3962));
XOR2_X1 i_3431 (.Z (n_3847), .A (n_2515), .B (n_3850));
XOR2_X1 i_3430 (.Z (n_2537), .A (n_2535), .B (n_3847));
AOI21_X1 i_3429 (.ZN (n_3846), .A (n_2415), .B1 (n_2414), .B2 (n_3982));
INV_X1 i_3428 (.ZN (n_2418), .A (n_3846));
AOI21_X1 i_3427 (.ZN (n_3845), .A (n_2405), .B1 (n_2404), .B2 (n_3958));
INV_X1 i_3426 (.ZN (n_3844), .A (n_3845));
XNOR2_X1 i_3425 (.ZN (n_2542), .A (n_2540), .B (n_3845));
AOI21_X1 i_3424 (.ZN (n_3843), .A (n_2420), .B1 (n_2419), .B2 (n_3957));
INV_X1 i_3423 (.ZN (n_2423), .A (n_3843));
AOI21_X1 i_3422 (.ZN (n_3842), .A (n_2430), .B1 (n_2429), .B2 (n_3952));
INV_X1 i_3421 (.ZN (n_2433), .A (n_3842));
AOI22_X1 i_3420 (.ZN (n_3841), .A1 (inputB[10]), .A2 (inputA[14]), .B1 (inputB[11]), .B2 (inputA[13]));
NAND3_X1 i_3419 (.ZN (n_3840), .A1 (inputB[11]), .A2 (inputA[14]), .A3 (n_4032));
INV_X1 i_3418 (.ZN (n_3839), .A (n_3840));
NOR2_X1 i_3417 (.ZN (n_3838), .A1 (n_3841), .A2 (n_3839));
NAND2_X1 i_3416 (.ZN (n_3837), .A1 (inputB[12]), .A2 (inputA[12]));
XNOR2_X1 i_3415 (.ZN (n_3836), .A (n_3838), .B (n_3837));
XOR2_X1 i_3414 (.Z (n_3833), .A (n_2525), .B (n_3836));
XOR2_X1 i_3413 (.Z (n_2552), .A (n_2550), .B (n_3833));
AOI21_X1 i_3412 (.ZN (n_3832), .A (n_2425), .B1 (n_2424), .B2 (n_3937));
INV_X1 i_3411 (.ZN (n_3831), .A (n_3832));
XNOR2_X1 i_3410 (.ZN (n_2562), .A (n_2560), .B (n_3832));
AOI21_X1 i_3409 (.ZN (n_3830), .A (n_2435), .B1 (n_2434), .B2 (n_3936));
INV_X1 i_3408 (.ZN (n_2438), .A (n_3830));
AOI21_X1 i_3407 (.ZN (n_3829), .A (n_2440), .B1 (n_2439), .B2 (n_3933));
INV_X1 i_3406 (.ZN (n_2443), .A (n_3829));
NAND3_X1 i_3405 (.ZN (n_3826), .A1 (inputB[2]), .A2 (inputA[23]), .A3 (n_4146));
AOI22_X1 i_3404 (.ZN (n_3825), .A1 (inputB[1]), .A2 (inputA[23]), .B1 (inputB[2]), .B2 (inputA[22]));
INV_X1 i_3403 (.ZN (n_3824), .A (n_3825));
NAND2_X1 i_3402 (.ZN (n_3823), .A1 (n_3826), .A2 (n_3824));
NAND2_X1 i_3401 (.ZN (n_3822), .A1 (inputB[3]), .A2 (inputA[21]));
XOR2_X1 i_3400 (.Z (n_3821), .A (n_3823), .B (n_3822));
XOR2_X1 i_3399 (.Z (n_3820), .A (n_2520), .B (n_3821));
XOR2_X1 i_3398 (.Z (n_3819), .A (n_2545), .B (n_3820));
XOR2_X1 i_3397 (.Z (n_3818), .A (n_2555), .B (n_3819));
XOR2_X1 i_3396 (.Z (n_3817), .A (n_2565), .B (n_3818));
XOR2_X1 i_3395 (.Z (n_2572), .A (n_2570), .B (n_3817));
AOI22_X1 i_3394 (.ZN (n_2491), .A1 (n_3995), .A2 (n_3922), .B1 (n_3916), .B2 (n_3912));
OAI21_X1 i_3393 (.ZN (n_2484), .A (n_3896), .B1 (n_3911), .B2 (n_3892));
OAI21_X1 i_3392 (.ZN (n_2470), .A (n_3886), .B1 (n_3888), .B2 (n_3884));
OAI21_X1 i_3391 (.ZN (n_2463), .A (n_3881), .B1 (n_3883), .B2 (n_3879));
OAI21_X1 i_3390 (.ZN (n_2449), .A (n_3874), .B1 (n_3878), .B2 (n_3872));
AOI21_X1 i_3389 (.ZN (n_3815), .A (n_2516), .B1 (n_2515), .B2 (n_3850));
INV_X1 i_3388 (.ZN (n_2519), .A (n_3815));
NOR2_X1 i_3387 (.ZN (n_3810), .A1 (n_3864), .A2 (n_3862));
AOI21_X1 i_3386 (.ZN (n_2505), .A (n_3810), .B1 (n_3866), .B2 (n_3865));
AND2_X1 i_3385 (.ZN (n_3806), .A1 (inputB[0]), .A2 (inputA[25]));
OAI21_X1 i_3384 (.ZN (n_3805), .A (n_3826), .B1 (n_3825), .B2 (n_3822));
NOR2_X1 i_3383 (.ZN (n_3800), .A1 (n_3806), .A2 (n_3805));
NAND2_X1 i_3382 (.ZN (n_3796), .A1 (n_3806), .A2 (n_3805));
OAI21_X1 i_3381 (.ZN (n_3795), .A (n_3796), .B1 (n_3806), .B2 (n_3805));
NAND2_X1 i_3380 (.ZN (n_3794), .A1 (inputB[1]), .A2 (inputA[24]));
XOR2_X1 i_3379 (.Z (n_2634), .A (n_3795), .B (n_3794));
AOI22_X1 i_3378 (.ZN (n_3790), .A1 (inputB[5]), .A2 (inputA[20]), .B1 (inputB[6]), .B2 (inputA[19]));
INV_X1 i_3377 (.ZN (n_3785), .A (n_3790));
NAND2_X1 i_3376 (.ZN (n_3784), .A1 (inputB[6]), .A2 (inputA[20]));
INV_X1 i_3375 (.ZN (n_3781), .A (n_3784));
NAND2_X1 i_3374 (.ZN (n_3780), .A1 (n_3917), .A2 (n_3781));
NAND2_X1 i_3373 (.ZN (n_3775), .A1 (n_3785), .A2 (n_3780));
NAND2_X1 i_3372 (.ZN (n_3770), .A1 (inputB[7]), .A2 (inputA[18]));
XOR2_X1 i_3371 (.Z (n_2621), .A (n_3775), .B (n_3770));
NAND2_X1 i_3370 (.ZN (n_3766), .A1 (inputB[9]), .A2 (inputA[16]));
INV_X1 i_3369 (.ZN (n_3765), .A (n_3766));
NAND2_X1 i_3368 (.ZN (n_3764), .A1 (n_3897), .A2 (n_3765));
OAI21_X1 i_3367 (.ZN (n_3760), .A (n_3764), .B1 (n_3897), .B2 (n_3765));
NAND2_X1 i_3365 (.ZN (n_3759), .A1 (inputB[10]), .A2 (inputA[15]));
XOR2_X1 i_3364 (.Z (n_2614), .A (n_3760), .B (n_3759));
AOI22_X1 i_3363 (.ZN (n_3756), .A1 (inputB[14]), .A2 (inputA[11]), .B1 (inputB[15]), .B2 (inputA[10]));
INV_X1 i_3361 (.ZN (n_3755), .A (n_3756));
NAND4_X1 i_3360 (.ZN (n_3750), .A1 (inputB[14]), .A2 (inputA[11]), .A3 (inputB[15]), .A4 (inputA[10]));
NAND2_X1 i_3359 (.ZN (n_3745), .A1 (n_3755), .A2 (n_3750));
NAND2_X1 i_3357 (.ZN (n_3744), .A1 (inputB[16]), .A2 (inputA[9]));
XOR2_X1 i_3356 (.Z (n_2600), .A (n_3745), .B (n_3744));
AND2_X1 i_3355 (.ZN (n_3740), .A1 (inputB[18]), .A2 (inputA[7]));
AOI21_X1 i_3353 (.ZN (n_3739), .A (n_3740), .B1 (inputB[17]), .B2 (inputA[8]));
INV_X1 i_3352 (.ZN (n_3735), .A (n_3739));
NAND3_X1 i_3351 (.ZN (n_3731), .A1 (inputB[17]), .A2 (inputA[8]), .A3 (n_3740));
NAND2_X1 i_3349 (.ZN (n_3730), .A1 (n_3735), .A2 (n_3731));
NAND2_X1 i_3348 (.ZN (n_3729), .A1 (inputB[19]), .A2 (inputA[6]));
XOR2_X1 i_3347 (.Z (n_2593), .A (n_3730), .B (n_3729));
AOI22_X1 i_3345 (.ZN (n_3725), .A1 (inputB[23]), .A2 (inputA[2]), .B1 (inputB[24]), .B2 (inputA[1]));
INV_X1 i_3344 (.ZN (n_3721), .A (n_3725));
NAND4_X1 i_3343 (.ZN (n_3720), .A1 (inputB[23]), .A2 (inputA[2]), .A3 (inputB[24]), .A4 (inputA[1]));
NAND2_X1 i_3341 (.ZN (n_3719), .A1 (n_3721), .A2 (n_3720));
NAND2_X1 i_3340 (.ZN (n_3718), .A1 (inputB[25]), .A2 (inputA[0]));
XOR2_X1 i_3339 (.Z (n_2579), .A (n_3719), .B (n_3718));
OAI21_X1 i_3337 (.ZN (n_3715), .A (n_3854), .B1 (n_3858), .B2 (n_3852));
XOR2_X1 i_3336 (.Z (n_2648), .A (n_2646), .B (n_3715));
AOI21_X1 i_3335 (.ZN (n_3714), .A (n_2531), .B1 (n_2530), .B2 (n_3851));
INV_X1 i_3333 (.ZN (n_2534), .A (n_3714));
AOI21_X1 i_3332 (.ZN (n_3713), .A (n_2526), .B1 (n_2525), .B2 (n_3836));
INV_X1 i_3331 (.ZN (n_2529), .A (n_3713));
AOI21_X1 i_3329 (.ZN (n_3712), .A (n_2511), .B1 (n_2510), .B2 (n_3868));
INV_X1 i_3328 (.ZN (n_3711), .A (n_3712));
XNOR2_X1 i_3327 (.ZN (n_2653), .A (n_2651), .B (n_3712));
AOI21_X1 i_3325 (.ZN (n_3709), .A (n_2541), .B1 (n_2540), .B2 (n_3844));
INV_X1 i_3324 (.ZN (n_2544), .A (n_3709));
AOI22_X1 i_3323 (.ZN (n_3708), .A1 (inputB[20]), .A2 (inputA[5]), .B1 (inputB[21]), .B2 (inputA[4]));
INV_X1 i_3321 (.ZN (n_3707), .A (n_3708));
AND2_X1 i_3320 (.ZN (n_3706), .A1 (inputB[21]), .A2 (inputA[5]));
NAND3_X1 i_3319 (.ZN (n_3705), .A1 (inputB[20]), .A2 (inputA[4]), .A3 (n_3706));
NAND2_X1 i_3317 (.ZN (n_3704), .A1 (n_3707), .A2 (n_3705));
NAND2_X1 i_3316 (.ZN (n_3701), .A1 (inputB[22]), .A2 (inputA[3]));
XOR2_X1 i_3315 (.Z (n_3700), .A (n_3704), .B (n_3701));
XOR2_X1 i_3313 (.Z (n_2668), .A (n_2666), .B (n_3700));
NAND2_X1 i_3312 (.ZN (n_3699), .A1 (inputB[12]), .A2 (inputA[14]));
INV_X1 i_3311 (.ZN (n_3698), .A (n_3699));
NAND3_X1 i_3309 (.ZN (n_3697), .A1 (inputB[11]), .A2 (inputA[13]), .A3 (n_3698));
AOI22_X1 i_3308 (.ZN (n_3696), .A1 (inputB[11]), .A2 (inputA[14]), .B1 (inputB[12]), .B2 (inputA[13]));
INV_X1 i_3307 (.ZN (n_3694), .A (n_3696));
NAND2_X1 i_3305 (.ZN (n_3693), .A1 (n_3697), .A2 (n_3694));
NAND2_X1 i_3304 (.ZN (n_3692), .A1 (inputB[13]), .A2 (inputA[12]));
XOR2_X1 i_3303 (.Z (n_3691), .A (n_3693), .B (n_3692));
XOR2_X1 i_3301 (.Z (n_2663), .A (n_2661), .B (n_3691));
AOI21_X1 i_3300 (.ZN (n_3690), .A (n_2546), .B1 (n_2545), .B2 (n_3820));
INV_X1 i_3299 (.ZN (n_2549), .A (n_3690));
AOI21_X1 i_3297 (.ZN (n_3688), .A (n_2521), .B1 (n_2520), .B2 (n_3821));
INV_X1 i_3296 (.ZN (n_3687), .A (n_3688));
XNOR2_X1 i_3295 (.ZN (n_2678), .A (n_2676), .B (n_3688));
AOI21_X1 i_3293 (.ZN (n_3686), .A (n_2551), .B1 (n_2550), .B2 (n_3833));
INV_X1 i_3292 (.ZN (n_2554), .A (n_3686));
AOI21_X1 i_3291 (.ZN (n_3685), .A (n_2536), .B1 (n_2535), .B2 (n_3847));
INV_X1 i_3290 (.ZN (n_3684), .A (n_3685));
XNOR2_X1 i_3289 (.ZN (n_2683), .A (n_2681), .B (n_3685));
AOI21_X1 i_3288 (.ZN (n_3683), .A (n_2561), .B1 (n_2560), .B2 (n_3831));
INV_X1 i_3287 (.ZN (n_2564), .A (n_3683));
NAND2_X1 i_3286 (.ZN (n_3680), .A1 (inputB[3]), .A2 (inputA[23]));
INV_X1 i_3285 (.ZN (n_3679), .A (n_3680));
NAND3_X1 i_3284 (.ZN (n_3678), .A1 (inputB[2]), .A2 (inputA[22]), .A3 (n_3679));
AOI22_X1 i_3283 (.ZN (n_3677), .A1 (inputB[2]), .A2 (inputA[23]), .B1 (inputB[3]), .B2 (inputA[22]));
INV_X1 i_3282 (.ZN (n_3676), .A (n_3677));
NAND2_X1 i_3281 (.ZN (n_3675), .A1 (n_3678), .A2 (n_3676));
NAND2_X1 i_3280 (.ZN (n_3673), .A1 (inputB[4]), .A2 (inputA[21]));
XOR2_X1 i_3279 (.Z (n_3672), .A (n_3675), .B (n_3673));
XOR2_X1 i_3278 (.Z (n_3671), .A (n_2656), .B (n_3672));
XOR2_X1 i_3277 (.Z (n_2688), .A (n_2686), .B (n_3671));
AOI21_X1 i_3276 (.ZN (n_3670), .A (n_2566), .B1 (n_2565), .B2 (n_3818));
INV_X1 i_3275 (.ZN (n_2569), .A (n_3670));
AOI21_X1 i_3274 (.ZN (n_3669), .A (n_2556), .B1 (n_2555), .B2 (n_3819));
INV_X1 i_3273 (.ZN (n_3667), .A (n_3669));
XNOR2_X1 i_3272 (.ZN (n_2698), .A (n_2696), .B (n_3669));
AOI21_X1 i_3271 (.ZN (n_3666), .A (n_2571), .B1 (n_2570), .B2 (n_3817));
INV_X1 i_3270 (.ZN (n_2574), .A (n_3666));
OAI21_X1 i_3269 (.ZN (n_2629), .A (n_3678), .B1 (n_3677), .B2 (n_3673));
OAI21_X1 i_3268 (.ZN (n_2622), .A (n_3780), .B1 (n_3790), .B2 (n_3770));
OAI21_X1 i_3267 (.ZN (n_2608), .A (n_3697), .B1 (n_3696), .B2 (n_3692));
OAI21_X1 i_3266 (.ZN (n_2601), .A (n_3750), .B1 (n_3756), .B2 (n_3744));
OAI21_X1 i_3265 (.ZN (n_2587), .A (n_3705), .B1 (n_3708), .B2 (n_3701));
OAI21_X1 i_3264 (.ZN (n_2580), .A (n_3720), .B1 (n_3725), .B2 (n_3718));
AOI21_X1 i_3263 (.ZN (n_3665), .A (n_3841), .B1 (n_3840), .B2 (n_3837));
AOI21_X1 i_3262 (.ZN (n_3664), .A (n_2642), .B1 (n_2641), .B2 (n_3665));
INV_X1 i_3261 (.ZN (n_2645), .A (n_3664));
OAI21_X1 i_3260 (.ZN (n_2635), .A (n_3796), .B1 (n_3800), .B2 (n_3794));
NAND2_X1 i_3259 (.ZN (n_3663), .A1 (inputB[4]), .A2 (inputA[22]));
INV_X1 i_3258 (.ZN (n_3662), .A (n_3663));
NAND2_X1 i_3257 (.ZN (n_3659), .A1 (n_3680), .A2 (n_3663));
AOI22_X1 i_3256 (.ZN (n_3658), .A1 (n_3679), .A2 (n_3662), .B1 (n_3680), .B2 (n_3663));
AND2_X1 i_3255 (.ZN (n_3657), .A1 (inputB[5]), .A2 (inputA[21]));
XOR2_X1 i_3254 (.Z (n_2764), .A (n_3658), .B (n_3657));
NAND2_X1 i_3253 (.ZN (n_3656), .A1 (inputB[7]), .A2 (inputA[19]));
INV_X1 i_3252 (.ZN (n_3655), .A (n_3656));
NAND2_X1 i_3251 (.ZN (n_3654), .A1 (n_3781), .A2 (n_3655));
NAND2_X1 i_3250 (.ZN (n_3652), .A1 (n_3784), .A2 (n_3656));
AND2_X1 i_3249 (.ZN (n_3651), .A1 (n_3654), .A2 (n_3652));
AND2_X1 i_3248 (.ZN (n_3650), .A1 (inputB[8]), .A2 (inputA[18]));
XOR2_X1 i_3247 (.Z (n_2757), .A (n_3651), .B (n_3650));
NAND2_X1 i_3246 (.ZN (n_3648), .A1 (inputB[13]), .A2 (inputA[13]));
INV_X1 i_3245 (.ZN (n_3647), .A (n_3648));
NAND2_X1 i_3244 (.ZN (n_3644), .A1 (n_3698), .A2 (n_3647));
NAND2_X1 i_3243 (.ZN (n_3643), .A1 (n_3699), .A2 (n_3648));
AND2_X1 i_3242 (.ZN (n_3639), .A1 (n_3644), .A2 (n_3643));
AND2_X1 i_3241 (.ZN (n_3638), .A1 (inputB[14]), .A2 (inputA[12]));
XOR2_X1 i_3240 (.Z (n_2743), .A (n_3639), .B (n_3638));
AND2_X1 i_3239 (.ZN (n_3637), .A1 (inputB[16]), .A2 (inputA[10]));
AOI21_X1 i_3238 (.ZN (n_3633), .A (n_3637), .B1 (inputB[15]), .B2 (inputA[11]));
INV_X1 i_3237 (.ZN (n_3628), .A (n_3633));
NAND3_X1 i_3236 (.ZN (n_3627), .A1 (inputB[15]), .A2 (inputA[11]), .A3 (n_3637));
NAND2_X1 i_3235 (.ZN (n_3623), .A1 (n_3628), .A2 (n_3627));
NAND2_X1 i_3234 (.ZN (n_3619), .A1 (inputB[17]), .A2 (inputA[9]));
XOR2_X1 i_3233 (.Z (n_2736), .A (n_3623), .B (n_3619));
AOI21_X1 i_3232 (.ZN (n_3618), .A (n_3706), .B1 (inputB[22]), .B2 (inputA[4]));
INV_X1 i_3231 (.ZN (n_3613), .A (n_3618));
NAND3_X1 i_3230 (.ZN (n_3608), .A1 (inputB[22]), .A2 (inputA[4]), .A3 (n_3706));
NAND2_X1 i_3229 (.ZN (n_3603), .A1 (n_3613), .A2 (n_3608));
NAND2_X1 i_3228 (.ZN (n_3598), .A1 (inputB[23]), .A2 (inputA[3]));
XOR2_X1 i_3227 (.Z (n_2722), .A (n_3603), .B (n_3598));
AND2_X1 i_3226 (.ZN (n_3597), .A1 (inputB[25]), .A2 (inputA[1]));
AOI21_X1 i_3225 (.ZN (n_3593), .A (n_3597), .B1 (inputB[24]), .B2 (inputA[2]));
INV_X1 i_3224 (.ZN (n_3588), .A (n_3593));
NAND3_X1 i_3223 (.ZN (n_3587), .A1 (inputB[24]), .A2 (inputA[2]), .A3 (n_3597));
NAND2_X1 i_3222 (.ZN (n_3584), .A1 (n_3588), .A2 (n_3587));
NAND2_X1 i_3221 (.ZN (n_3583), .A1 (inputB[26]), .A2 (inputA[0]));
XOR2_X1 i_3220 (.Z (n_2715), .A (n_3584), .B (n_3583));
AOI21_X1 i_3219 (.ZN (n_3578), .A (n_2647), .B1 (n_2646), .B2 (n_3715));
INV_X1 i_3218 (.ZN (n_3573), .A (n_3578));
XNOR2_X1 i_3217 (.ZN (n_2788), .A (n_2786), .B (n_3578));
OAI21_X1 i_3216 (.ZN (n_3568), .A (n_3731), .B1 (n_3739), .B2 (n_3729));
XOR2_X1 i_3215 (.Z (n_2783), .A (n_2781), .B (n_3568));
AOI21_X1 i_3213 (.ZN (n_3563), .A (n_2667), .B1 (n_2666), .B2 (n_3700));
INV_X1 i_3212 (.ZN (n_2670), .A (n_3563));
AOI21_X1 i_3211 (.ZN (n_3559), .A (n_2662), .B1 (n_2661), .B2 (n_3691));
INV_X1 i_3209 (.ZN (n_2665), .A (n_3559));
AOI22_X1 i_3208 (.ZN (n_3558), .A1 (inputB[0]), .A2 (inputA[26]), .B1 (inputB[1]), .B2 (inputA[25]));
INV_X1 i_3207 (.ZN (n_3557), .A (n_3558));
NAND3_X1 i_3205 (.ZN (n_3554), .A1 (inputB[1]), .A2 (inputA[26]), .A3 (n_3806));
NAND2_X1 i_3204 (.ZN (n_3553), .A1 (n_3557), .A2 (n_3554));
NAND2_X1 i_3203 (.ZN (n_3552), .A1 (inputB[2]), .A2 (inputA[24]));
XOR2_X1 i_3201 (.Z (n_3551), .A (n_3553), .B (n_3552));
XOR2_X1 i_3200 (.Z (n_2793), .A (n_2791), .B (n_3551));
AOI21_X1 i_3199 (.ZN (n_3548), .A (n_2677), .B1 (n_2676), .B2 (n_3687));
INV_X1 i_3197 (.ZN (n_2680), .A (n_3548));
AOI21_X1 i_3196 (.ZN (n_3547), .A (n_2652), .B1 (n_2651), .B2 (n_3711));
INV_X1 i_3195 (.ZN (n_3546), .A (n_3547));
XNOR2_X1 i_3193 (.ZN (n_2808), .A (n_2806), .B (n_3547));
NAND2_X1 i_3192 (.ZN (n_3545), .A1 (inputB[19]), .A2 (inputA[8]));
INV_X1 i_3191 (.ZN (n_3544), .A (n_3545));
NAND2_X1 i_3189 (.ZN (n_3543), .A1 (n_3740), .A2 (n_3544));
AOI22_X1 i_3188 (.ZN (n_3541), .A1 (inputB[18]), .A2 (inputA[8]), .B1 (inputB[19]), .B2 (inputA[7]));
INV_X1 i_3187 (.ZN (n_3540), .A (n_3541));
NAND2_X1 i_3185 (.ZN (n_3539), .A1 (n_3543), .A2 (n_3540));
NAND2_X1 i_3184 (.ZN (n_3538), .A1 (inputB[20]), .A2 (inputA[6]));
XOR2_X1 i_3183 (.Z (n_3537), .A (n_3539), .B (n_3538));
XOR2_X1 i_3181 (.Z (n_2803), .A (n_2801), .B (n_3537));
AOI21_X1 i_3180 (.ZN (n_3535), .A (n_2682), .B1 (n_2681), .B2 (n_3684));
INV_X1 i_3179 (.ZN (n_2685), .A (n_3535));
AOI21_X1 i_3177 (.ZN (n_3534), .A (n_2657), .B1 (n_2656), .B2 (n_3672));
INV_X1 i_3176 (.ZN (n_3533), .A (n_3534));
XNOR2_X1 i_3175 (.ZN (n_2818), .A (n_2816), .B (n_3534));
AOI21_X1 i_3173 (.ZN (n_3532), .A (n_2687), .B1 (n_2686), .B2 (n_3671));
INV_X1 i_3172 (.ZN (n_2690), .A (n_3532));
XOR2_X1 i_3171 (.Z (n_3531), .A (n_2641), .B (n_3665));
AOI21_X1 i_3169 (.ZN (n_3530), .A (n_2672), .B1 (n_2671), .B2 (n_3531));
INV_X1 i_3168 (.ZN (n_3527), .A (n_3530));
XNOR2_X1 i_3167 (.ZN (n_2823), .A (n_2821), .B (n_3530));
NAND2_X1 i_3165 (.ZN (n_3526), .A1 (inputB[10]), .A2 (inputA[17]));
INV_X1 i_3164 (.ZN (n_3525), .A (n_3526));
NAND2_X1 i_3163 (.ZN (n_3524), .A1 (n_3765), .A2 (n_3525));
AOI22_X1 i_3161 (.ZN (n_3523), .A1 (inputB[9]), .A2 (inputA[17]), .B1 (inputB[10]), .B2 (inputA[16]));
INV_X1 i_3160 (.ZN (n_3522), .A (n_3523));
NAND2_X1 i_3159 (.ZN (n_3520), .A1 (n_3524), .A2 (n_3522));
NAND2_X1 i_3157 (.ZN (n_3519), .A1 (inputB[11]), .A2 (inputA[15]));
XOR2_X1 i_3156 (.Z (n_3518), .A (n_3520), .B (n_3519));
XOR2_X1 i_3155 (.Z (n_3517), .A (n_2796), .B (n_3518));
XOR2_X1 i_3153 (.Z (n_2828), .A (n_2826), .B (n_3517));
AOI21_X1 i_3152 (.ZN (n_3516), .A (n_2697), .B1 (n_2696), .B2 (n_3667));
INV_X1 i_3151 (.ZN (n_2700), .A (n_3516));
XOR2_X1 i_3149 (.Z (n_3514), .A (n_2671), .B (n_3531));
AOI21_X1 i_3148 (.ZN (n_3513), .A (n_2692), .B1 (n_2691), .B2 (n_3514));
INV_X1 i_3147 (.ZN (n_3512), .A (n_3513));
XNOR2_X1 i_3145 (.ZN (n_2838), .A (n_2836), .B (n_3513));
XOR2_X1 i_3144 (.Z (n_3511), .A (n_2691), .B (n_3514));
AOI21_X1 i_3143 (.ZN (n_3510), .A (n_2702), .B1 (n_2701), .B2 (n_3511));
INV_X1 i_3142 (.ZN (n_2705), .A (n_3510));
XOR2_X1 i_3141 (.Z (n_3509), .A (n_2701), .B (n_3511));
AOI21_X1 i_3140 (.ZN (n_3506), .A (n_2707), .B1 (n_2706), .B2 (n_3509));
INV_X1 i_3139 (.ZN (n_2710), .A (n_3506));
AOI22_X1 i_3138 (.ZN (n_3505), .A1 (n_3902), .A2 (n_3766), .B1 (n_3764), .B2 (n_3759));
XOR2_X1 i_3137 (.Z (n_3504), .A (n_2776), .B (n_3505));
XOR2_X1 i_3136 (.Z (n_3503), .A (n_2811), .B (n_3504));
XOR2_X1 i_3135 (.Z (n_3502), .A (n_2831), .B (n_3503));
XOR2_X1 i_3134 (.Z (n_3501), .A (n_2841), .B (n_3502));
XOR2_X1 i_3133 (.Z (n_2848), .A (n_2846), .B (n_3501));
NAND2_X1 i_3132 (.ZN (n_3499), .A1 (n_3652), .A2 (n_3650));
NAND2_X1 i_3131 (.ZN (n_2758), .A1 (n_3654), .A2 (n_3499));
OAI21_X1 i_3130 (.ZN (n_2751), .A (n_3524), .B1 (n_3523), .B2 (n_3519));
OAI21_X1 i_3129 (.ZN (n_2737), .A (n_3627), .B1 (n_3633), .B2 (n_3619));
OAI21_X1 i_3128 (.ZN (n_2730), .A (n_3543), .B1 (n_3541), .B2 (n_3538));
OAI21_X1 i_3127 (.ZN (n_2716), .A (n_3587), .B1 (n_3593), .B2 (n_3583));
AOI21_X1 i_3126 (.ZN (n_3498), .A (n_2782), .B1 (n_2781), .B2 (n_3568));
INV_X1 i_3125 (.ZN (n_2785), .A (n_3498));
AND2_X1 i_3124 (.ZN (n_3497), .A1 (inputB[2]), .A2 (inputA[26]));
NAND3_X1 i_3123 (.ZN (n_3496), .A1 (inputB[1]), .A2 (inputA[25]), .A3 (n_3497));
AOI22_X1 i_3122 (.ZN (n_3495), .A1 (inputB[1]), .A2 (inputA[26]), .B1 (inputB[2]), .B2 (inputA[25]));
INV_X1 i_3121 (.ZN (n_3493), .A (n_3495));
NAND2_X1 i_3120 (.ZN (n_3492), .A1 (n_3496), .A2 (n_3493));
NAND2_X1 i_3119 (.ZN (n_3491), .A1 (inputB[3]), .A2 (inputA[24]));
XOR2_X1 i_3118 (.Z (n_2911), .A (n_3492), .B (n_3491));
AOI22_X1 i_3117 (.ZN (n_3490), .A1 (inputB[4]), .A2 (inputA[23]), .B1 (inputB[5]), .B2 (inputA[22]));
INV_X1 i_3116 (.ZN (n_3489), .A (n_3490));
NAND2_X1 i_3115 (.ZN (n_3488), .A1 (inputB[5]), .A2 (inputA[23]));
INV_X1 i_3114 (.ZN (n_3485), .A (n_3488));
NAND2_X1 i_3113 (.ZN (n_3484), .A1 (n_3662), .A2 (n_3485));
NAND2_X1 i_3112 (.ZN (n_3483), .A1 (n_3489), .A2 (n_3484));
NAND2_X1 i_3111 (.ZN (n_3482), .A1 (inputB[6]), .A2 (inputA[21]));
XOR2_X1 i_3110 (.Z (n_2904), .A (n_3483), .B (n_3482));
NAND2_X1 i_3109 (.ZN (n_3481), .A1 (inputB[11]), .A2 (inputA[16]));
INV_X1 i_3108 (.ZN (n_3480), .A (n_3481));
NAND2_X1 i_3107 (.ZN (n_3479), .A1 (n_3525), .A2 (n_3480));
OAI21_X1 i_3106 (.ZN (n_3478), .A (n_3479), .B1 (n_3525), .B2 (n_3480));
NAND2_X1 i_3105 (.ZN (n_3476), .A1 (inputB[12]), .A2 (inputA[15]));
XOR2_X1 i_3104 (.Z (n_2890), .A (n_3478), .B (n_3476));
AOI22_X1 i_3103 (.ZN (n_3472), .A1 (inputB[13]), .A2 (inputA[14]), .B1 (inputB[14]), .B2 (inputA[13]));
INV_X1 i_3102 (.ZN (n_3467), .A (n_3472));
NAND2_X1 i_3101 (.ZN (n_3466), .A1 (inputB[14]), .A2 (inputA[14]));
INV_X1 i_3100 (.ZN (n_3462), .A (n_3466));
NAND2_X1 i_3099 (.ZN (n_3458), .A1 (n_3647), .A2 (n_3462));
NAND2_X1 i_3098 (.ZN (n_3457), .A1 (n_3467), .A2 (n_3458));
NAND2_X1 i_3097 (.ZN (n_3453), .A1 (inputB[15]), .A2 (inputA[12]));
XOR2_X1 i_3096 (.Z (n_2883), .A (n_3457), .B (n_3453));
NAND2_X1 i_3095 (.ZN (n_3452), .A1 (inputB[20]), .A2 (inputA[7]));
INV_X1 i_3094 (.ZN (n_3447), .A (n_3452));
NAND2_X1 i_3093 (.ZN (n_3443), .A1 (n_3544), .A2 (n_3447));
OAI21_X1 i_3092 (.ZN (n_3442), .A (n_3443), .B1 (n_3544), .B2 (n_3447));
NAND2_X1 i_3091 (.ZN (n_3441), .A1 (inputB[21]), .A2 (inputA[6]));
XOR2_X1 i_3090 (.Z (n_2869), .A (n_3442), .B (n_3441));
AOI22_X1 i_3089 (.ZN (n_3437), .A1 (inputB[22]), .A2 (inputA[5]), .B1 (inputB[23]), .B2 (inputA[4]));
INV_X1 i_3088 (.ZN (n_3433), .A (n_3437));
NAND4_X1 i_3087 (.ZN (n_3432), .A1 (inputB[22]), .A2 (inputA[5]), .A3 (inputB[23]), .A4 (inputA[4]));
NAND2_X1 i_3086 (.ZN (n_3431), .A1 (n_3433), .A2 (n_3432));
NAND2_X1 i_3085 (.ZN (n_3427), .A1 (inputB[24]), .A2 (inputA[3]));
XOR2_X1 i_3084 (.Z (n_2862), .A (n_3431), .B (n_3427));
AOI21_X1 i_3083 (.ZN (n_3422), .A (n_2787), .B1 (n_2786), .B2 (n_3573));
INV_X1 i_3082 (.ZN (n_2790), .A (n_3422));
OAI21_X1 i_3081 (.ZN (n_3417), .A (n_3608), .B1 (n_3618), .B2 (n_3598));
XOR2_X1 i_3080 (.Z (n_2931), .A (n_2929), .B (n_3417));
OAI21_X1 i_3079 (.ZN (n_3413), .A (n_3554), .B1 (n_3558), .B2 (n_3552));
INV_X1 i_3078 (.ZN (n_3412), .A (n_3413));
AOI22_X1 i_3077 (.ZN (n_3411), .A1 (n_3679), .A2 (n_3662), .B1 (n_3659), .B2 (n_3657));
NOR2_X1 i_3076 (.ZN (n_3407), .A1 (n_3412), .A2 (n_3411));
AOI21_X1 i_3075 (.ZN (n_3406), .A (n_3407), .B1 (n_3412), .B2 (n_3411));
AND2_X1 i_3074 (.ZN (n_3403), .A1 (inputB[0]), .A2 (inputA[27]));
XOR2_X1 i_3073 (.Z (n_2918), .A (n_3406), .B (n_3403));
AOI21_X1 i_3072 (.ZN (n_3402), .A (n_2802), .B1 (n_2801), .B2 (n_3537));
INV_X1 i_3071 (.ZN (n_2805), .A (n_3402));
AOI21_X1 i_3070 (.ZN (n_3397), .A (n_2792), .B1 (n_2791), .B2 (n_3551));
INV_X1 i_3069 (.ZN (n_2795), .A (n_3397));
AOI21_X1 i_3068 (.ZN (n_3396), .A (n_2807), .B1 (n_2806), .B2 (n_3546));
INV_X1 i_3066 (.ZN (n_2810), .A (n_3396));
AOI21_X1 i_3065 (.ZN (n_3392), .A (n_2817), .B1 (n_2816), .B2 (n_3533));
INV_X1 i_3064 (.ZN (n_2820), .A (n_3392));
AOI21_X1 i_3062 (.ZN (n_3388), .A (n_2812), .B1 (n_2811), .B2 (n_3504));
INV_X1 i_3061 (.ZN (n_2815), .A (n_3388));
AOI22_X1 i_3060 (.ZN (n_3387), .A1 (inputB[16]), .A2 (inputA[11]), .B1 (inputB[17]), .B2 (inputA[10]));
INV_X1 i_3058 (.ZN (n_3386), .A (n_3387));
NAND3_X1 i_3057 (.ZN (n_3385), .A1 (inputB[17]), .A2 (inputA[11]), .A3 (n_3637));
NAND2_X1 i_3056 (.ZN (n_3384), .A1 (n_3386), .A2 (n_3385));
NAND2_X1 i_3054 (.ZN (n_3382), .A1 (inputB[18]), .A2 (inputA[9]));
XOR2_X1 i_3053 (.Z (n_3381), .A (n_3384), .B (n_3382));
XOR2_X1 i_3052 (.Z (n_2946), .A (n_2944), .B (n_3381));
NAND3_X1 i_3050 (.ZN (n_3380), .A1 (inputB[8]), .A2 (inputA[20]), .A3 (n_3655));
AOI22_X1 i_3049 (.ZN (n_3379), .A1 (inputB[7]), .A2 (inputA[20]), .B1 (inputB[8]), .B2 (inputA[19]));
INV_X1 i_3048 (.ZN (n_3378), .A (n_3379));
NAND2_X1 i_3046 (.ZN (n_3377), .A1 (n_3380), .A2 (n_3378));
NAND2_X1 i_3045 (.ZN (n_3376), .A1 (inputB[9]), .A2 (inputA[18]));
XOR2_X1 i_3044 (.Z (n_3375), .A (n_3377), .B (n_3376));
XOR2_X1 i_3042 (.Z (n_2941), .A (n_2939), .B (n_3375));
AOI21_X1 i_3041 (.ZN (n_3374), .A (n_2797), .B1 (n_2796), .B2 (n_3518));
INV_X1 i_3040 (.ZN (n_3373), .A (n_3374));
XNOR2_X1 i_3038 (.ZN (n_2961), .A (n_2959), .B (n_3374));
NAND2_X1 i_3037 (.ZN (n_3372), .A1 (n_3643), .A2 (n_3638));
NAND2_X1 i_3036 (.ZN (n_3371), .A1 (n_3644), .A2 (n_3372));
XOR2_X1 i_3034 (.Z (n_3368), .A (n_2924), .B (n_3371));
XOR2_X1 i_3033 (.Z (n_2956), .A (n_2954), .B (n_3368));
AOI21_X1 i_3032 (.ZN (n_3367), .A (n_2777), .B1 (n_2776), .B2 (n_3505));
INV_X1 i_3030 (.ZN (n_3366), .A (n_3367));
XNOR2_X1 i_3029 (.ZN (n_3365), .A (n_2934), .B (n_3367));
XOR2_X1 i_3028 (.Z (n_2966), .A (n_2964), .B (n_3365));
NAND2_X1 i_3026 (.ZN (n_3364), .A1 (inputB[26]), .A2 (inputA[2]));
INV_X1 i_3025 (.ZN (n_3361), .A (n_3364));
NAND2_X1 i_3024 (.ZN (n_3360), .A1 (n_3597), .A2 (n_3361));
AOI22_X1 i_3022 (.ZN (n_3359), .A1 (inputB[25]), .A2 (inputA[2]), .B1 (inputB[26]), .B2 (inputA[1]));
INV_X1 i_3021 (.ZN (n_3358), .A (n_3359));
NAND2_X1 i_3020 (.ZN (n_3357), .A1 (n_3360), .A2 (n_3358));
NAND2_X1 i_3018 (.ZN (n_3356), .A1 (inputB[27]), .A2 (inputA[0]));
XOR2_X1 i_3017 (.Z (n_3355), .A (n_3357), .B (n_3356));
XOR2_X1 i_3016 (.Z (n_3354), .A (n_2949), .B (n_3355));
XOR2_X1 i_3014 (.Z (n_2971), .A (n_2969), .B (n_3354));
AOI21_X1 i_3013 (.ZN (n_3353), .A (n_2822), .B1 (n_2821), .B2 (n_3527));
INV_X1 i_3012 (.ZN (n_3352), .A (n_3353));
XNOR2_X1 i_3010 (.ZN (n_2976), .A (n_2974), .B (n_3353));
AOI21_X1 i_3009 (.ZN (n_3351), .A (n_2837), .B1 (n_2836), .B2 (n_3512));
INV_X1 i_3008 (.ZN (n_2840), .A (n_3351));
AOI21_X1 i_3006 (.ZN (n_3350), .A (n_2832), .B1 (n_2831), .B2 (n_3503));
INV_X1 i_3005 (.ZN (n_3347), .A (n_3350));
XNOR2_X1 i_3004 (.ZN (n_2986), .A (n_2984), .B (n_3350));
AOI21_X1 i_3002 (.ZN (n_3346), .A (n_2842), .B1 (n_2841), .B2 (n_3502));
INV_X1 i_3001 (.ZN (n_2845), .A (n_3346));
AOI21_X1 i_3000 (.ZN (n_3345), .A (n_2847), .B1 (n_2846), .B2 (n_3501));
INV_X1 i_2998 (.ZN (n_2850), .A (n_3345));
AOI21_X1 i_2997 (.ZN (n_3344), .A (n_2827), .B1 (n_2826), .B2 (n_3517));
INV_X1 i_2996 (.ZN (n_3343), .A (n_3344));
XNOR2_X1 i_2995 (.ZN (n_3340), .A (n_2979), .B (n_3344));
XOR2_X1 i_2994 (.Z (n_3339), .A (n_2989), .B (n_3340));
XOR2_X1 i_2993 (.Z (n_2996), .A (n_2994), .B (n_3339));
OAI21_X1 i_2992 (.ZN (n_2905), .A (n_3484), .B1 (n_3490), .B2 (n_3482));
OAI21_X1 i_2991 (.ZN (n_2898), .A (n_3380), .B1 (n_3379), .B2 (n_3376));
OAI21_X1 i_2990 (.ZN (n_2884), .A (n_3458), .B1 (n_3472), .B2 (n_3453));
OAI21_X1 i_2989 (.ZN (n_2877), .A (n_3385), .B1 (n_3387), .B2 (n_3382));
OAI21_X1 i_2988 (.ZN (n_2863), .A (n_3432), .B1 (n_3437), .B2 (n_3427));
OAI21_X1 i_2987 (.ZN (n_2856), .A (n_3360), .B1 (n_3359), .B2 (n_3356));
AOI21_X1 i_2986 (.ZN (n_3338), .A (n_2925), .B1 (n_2924), .B2 (n_3371));
INV_X1 i_2985 (.ZN (n_2928), .A (n_3338));
NOR2_X1 i_2984 (.ZN (n_3337), .A1 (n_3407), .A2 (n_3403));
AOI21_X1 i_2983 (.ZN (n_2919), .A (n_3337), .B1 (n_3412), .B2 (n_3411));
NAND3_X1 i_2982 (.ZN (n_3336), .A1 (inputB[3]), .A2 (inputA[25]), .A3 (n_3497));
INV_X1 i_2981 (.ZN (n_3335), .A (n_3336));
AOI21_X1 i_2980 (.ZN (n_3334), .A (n_3497), .B1 (inputB[3]), .B2 (inputA[25]));
NOR2_X1 i_2979 (.ZN (n_3333), .A1 (n_3335), .A2 (n_3334));
NAND2_X1 i_2978 (.ZN (n_3332), .A1 (inputB[4]), .A2 (inputA[24]));
XNOR2_X1 i_2977 (.ZN (n_3059), .A (n_3333), .B (n_3332));
NAND2_X1 i_2976 (.ZN (n_3331), .A1 (inputB[6]), .A2 (inputA[22]));
INV_X1 i_2975 (.ZN (n_3330), .A (n_3331));
NAND2_X1 i_2974 (.ZN (n_3329), .A1 (n_3485), .A2 (n_3330));
OAI21_X1 i_2973 (.ZN (n_3326), .A (n_3329), .B1 (n_3485), .B2 (n_3330));
NAND2_X1 i_2972 (.ZN (n_3325), .A1 (inputB[7]), .A2 (inputA[21]));
XOR2_X1 i_2971 (.Z (n_3052), .A (n_3326), .B (n_3325));
AOI22_X1 i_2970 (.ZN (n_3324), .A1 (inputB[11]), .A2 (inputA[17]), .B1 (inputB[12]), .B2 (inputA[16]));
INV_X1 i_2969 (.ZN (n_3323), .A (n_3324));
AND2_X1 i_2968 (.ZN (n_3322), .A1 (inputB[12]), .A2 (inputA[17]));
NAND2_X1 i_2967 (.ZN (n_3319), .A1 (n_3480), .A2 (n_3322));
NAND2_X1 i_2966 (.ZN (n_3318), .A1 (n_3323), .A2 (n_3319));
NAND2_X1 i_2965 (.ZN (n_3317), .A1 (inputB[13]), .A2 (inputA[15]));
XOR2_X1 i_2964 (.Z (n_3038), .A (n_3318), .B (n_3317));
NAND2_X1 i_2963 (.ZN (n_3316), .A1 (inputB[15]), .A2 (inputA[13]));
INV_X1 i_2962 (.ZN (n_3315), .A (n_3316));
NAND2_X1 i_2961 (.ZN (n_3314), .A1 (n_3462), .A2 (n_3315));
OAI21_X1 i_2960 (.ZN (n_3313), .A (n_3314), .B1 (n_3462), .B2 (n_3315));
NAND2_X1 i_2959 (.ZN (n_3312), .A1 (inputB[16]), .A2 (inputA[12]));
XOR2_X1 i_2958 (.Z (n_3031), .A (n_3313), .B (n_3312));
AOI22_X1 i_2957 (.ZN (n_3311), .A1 (inputB[20]), .A2 (inputA[8]), .B1 (inputB[21]), .B2 (inputA[7]));
INV_X1 i_2956 (.ZN (n_3307), .A (n_3311));
AND2_X1 i_2955 (.ZN (n_3302), .A1 (inputB[21]), .A2 (inputA[8]));
NAND2_X1 i_2954 (.ZN (n_3301), .A1 (n_3447), .A2 (n_3302));
NAND2_X1 i_2953 (.ZN (n_3298), .A1 (n_3307), .A2 (n_3301));
NAND2_X1 i_2952 (.ZN (n_3297), .A1 (inputB[22]), .A2 (inputA[6]));
XOR2_X1 i_2951 (.Z (n_3017), .A (n_3298), .B (n_3297));
AND2_X1 i_2950 (.ZN (n_3293), .A1 (inputB[24]), .A2 (inputA[4]));
AOI21_X1 i_2949 (.ZN (n_3292), .A (n_3293), .B1 (inputB[23]), .B2 (inputA[5]));
INV_X1 i_2948 (.ZN (n_3287), .A (n_3292));
NAND3_X1 i_2947 (.ZN (n_3282), .A1 (inputB[23]), .A2 (inputA[5]), .A3 (n_3293));
NAND2_X1 i_2946 (.ZN (n_3281), .A1 (n_3287), .A2 (n_3282));
NAND2_X1 i_2945 (.ZN (n_3277), .A1 (inputB[25]), .A2 (inputA[3]));
XOR2_X1 i_2944 (.Z (n_3010), .A (n_3281), .B (n_3277));
AOI21_X1 i_2943 (.ZN (n_3276), .A (n_2935), .B1 (n_2934), .B2 (n_3366));
INV_X1 i_2942 (.ZN (n_2938), .A (n_3276));
AOI21_X1 i_2941 (.ZN (n_3272), .A (n_2930), .B1 (n_2929), .B2 (n_3417));
INV_X1 i_2940 (.ZN (n_3271), .A (n_3272));
XNOR2_X1 i_2939 (.ZN (n_3084), .A (n_3082), .B (n_3272));
AOI22_X1 i_2938 (.ZN (n_3267), .A1 (n_3526), .A2 (n_3481), .B1 (n_3479), .B2 (n_3476));
XOR2_X1 i_2937 (.Z (n_3074), .A (n_3072), .B (n_3267));
AOI21_X1 i_2936 (.ZN (n_3263), .A (n_2950), .B1 (n_2949), .B2 (n_3355));
INV_X1 i_2935 (.ZN (n_2953), .A (n_3263));
AOI21_X1 i_2934 (.ZN (n_3262), .A (n_2940), .B1 (n_2939), .B2 (n_3375));
INV_X1 i_2933 (.ZN (n_2943), .A (n_3262));
AND2_X1 i_2932 (.ZN (n_3258), .A1 (inputB[1]), .A2 (inputA[28]));
AOI22_X1 i_2931 (.ZN (n_3257), .A1 (inputB[0]), .A2 (inputA[28]), .B1 (inputB[1]), .B2 (inputA[27]));
AOI21_X1 i_2930 (.ZN (n_3252), .A (n_3257), .B1 (n_3403), .B2 (n_3258));
OAI21_X1 i_2929 (.ZN (n_3247), .A (n_3496), .B1 (n_3495), .B2 (n_3491));
XOR2_X1 i_2927 (.Z (n_3246), .A (n_3252), .B (n_3247));
XOR2_X1 i_2926 (.Z (n_3089), .A (n_3087), .B (n_3246));
AOI21_X1 i_2925 (.ZN (n_3242), .A (n_2955), .B1 (n_2954), .B2 (n_3368));
INV_X1 i_2923 (.ZN (n_2958), .A (n_3242));
NAND2_X1 i_2922 (.ZN (n_3238), .A1 (inputB[27]), .A2 (inputA[1]));
INV_X1 i_2921 (.ZN (n_3237), .A (n_3238));
NAND2_X1 i_2919 (.ZN (n_3236), .A1 (n_3361), .A2 (n_3237));
OAI21_X1 i_2918 (.ZN (n_3232), .A (n_3236), .B1 (n_3361), .B2 (n_3237));
NAND2_X1 i_2917 (.ZN (n_3227), .A1 (inputB[28]), .A2 (inputA[0]));
XOR2_X1 i_2915 (.Z (n_3223), .A (n_3232), .B (n_3227));
XOR2_X1 i_2914 (.Z (n_3104), .A (n_3102), .B (n_3223));
NAND2_X1 i_2913 (.ZN (n_3222), .A1 (inputB[9]), .A2 (inputA[20]));
INV_X1 i_2911 (.ZN (n_3221), .A (n_3222));
NAND3_X1 i_2910 (.ZN (n_3220), .A1 (inputB[8]), .A2 (inputA[19]), .A3 (n_3221));
INV_X1 i_2909 (.ZN (n_3218), .A (n_3220));
AOI22_X1 i_2907 (.ZN (n_3217), .A1 (inputB[8]), .A2 (inputA[20]), .B1 (inputB[9]), .B2 (inputA[19]));
NOR2_X1 i_2906 (.ZN (n_3216), .A1 (n_3218), .A2 (n_3217));
NAND2_X1 i_2905 (.ZN (n_3215), .A1 (inputB[10]), .A2 (inputA[18]));
XNOR2_X1 i_2903 (.ZN (n_3214), .A (n_3216), .B (n_3215));
XOR2_X1 i_2902 (.Z (n_3094), .A (n_3092), .B (n_3214));
AOI21_X1 i_2901 (.ZN (n_3213), .A (n_2965), .B1 (n_2964), .B2 (n_3365));
INV_X1 i_2899 (.ZN (n_2968), .A (n_3213));
AOI22_X1 i_2898 (.ZN (n_3211), .A1 (n_3545), .A2 (n_3452), .B1 (n_3443), .B2 (n_3441));
XOR2_X1 i_2897 (.Z (n_3210), .A (n_3077), .B (n_3211));
XOR2_X1 i_2895 (.Z (n_3109), .A (n_3107), .B (n_3210));
AOI21_X1 i_2894 (.ZN (n_3209), .A (n_2970), .B1 (n_2969), .B2 (n_3354));
INV_X1 i_2893 (.ZN (n_2973), .A (n_3209));
AOI21_X1 i_2891 (.ZN (n_3208), .A (n_2960), .B1 (n_2959), .B2 (n_3373));
INV_X1 i_2890 (.ZN (n_3207), .A (n_3208));
XNOR2_X1 i_2889 (.ZN (n_3119), .A (n_3117), .B (n_3208));
AOI21_X1 i_2887 (.ZN (n_3205), .A (n_2980), .B1 (n_2979), .B2 (n_3343));
INV_X1 i_2886 (.ZN (n_2983), .A (n_3205));
AOI21_X1 i_2885 (.ZN (n_3204), .A (n_2945), .B1 (n_2944), .B2 (n_3381));
INV_X1 i_2883 (.ZN (n_3203), .A (n_3204));
XNOR2_X1 i_2882 (.ZN (n_3202), .A (n_3112), .B (n_3204));
XOR2_X1 i_2881 (.Z (n_3129), .A (n_3127), .B (n_3202));
AOI21_X1 i_2879 (.ZN (n_3201), .A (n_2985), .B1 (n_2984), .B2 (n_3347));
INV_X1 i_2878 (.ZN (n_2988), .A (n_3201));
AOI22_X1 i_2877 (.ZN (n_3200), .A1 (inputB[17]), .A2 (inputA[11]), .B1 (inputB[18]), .B2 (inputA[10]));
NAND2_X1 i_2875 (.ZN (n_3197), .A1 (inputB[18]), .A2 (inputA[11]));
INV_X1 i_2874 (.ZN (n_3196), .A (n_3197));
NAND3_X1 i_2873 (.ZN (n_3195), .A1 (inputB[17]), .A2 (inputA[10]), .A3 (n_3196));
INV_X1 i_2871 (.ZN (n_3194), .A (n_3195));
NOR2_X1 i_2870 (.ZN (n_3193), .A1 (n_3200), .A2 (n_3194));
NAND2_X1 i_2869 (.ZN (n_3192), .A1 (inputB[19]), .A2 (inputA[9]));
XNOR2_X1 i_2867 (.ZN (n_3190), .A (n_3193), .B (n_3192));
XOR2_X1 i_2866 (.Z (n_3189), .A (n_3097), .B (n_3190));
XOR2_X1 i_2865 (.Z (n_3188), .A (n_3122), .B (n_3189));
XOR2_X1 i_2863 (.Z (n_3139), .A (n_3137), .B (n_3188));
AOI21_X1 i_2862 (.ZN (n_3187), .A (n_2990), .B1 (n_2989), .B2 (n_3340));
INV_X1 i_2861 (.ZN (n_2993), .A (n_3187));
AOI21_X1 i_2860 (.ZN (n_3186), .A (n_2995), .B1 (n_2994), .B2 (n_3339));
INV_X1 i_2859 (.ZN (n_2998), .A (n_3186));
AOI21_X1 i_2858 (.ZN (n_3184), .A (n_2975), .B1 (n_2974), .B2 (n_3352));
INV_X1 i_2857 (.ZN (n_3183), .A (n_3184));
XNOR2_X1 i_2856 (.ZN (n_3182), .A (n_3132), .B (n_3184));
XOR2_X1 i_2855 (.Z (n_3181), .A (n_3142), .B (n_3182));
XOR2_X1 i_2854 (.Z (n_3149), .A (n_3147), .B (n_3181));
OAI21_X1 i_2853 (.ZN (n_3060), .A (n_3336), .B1 (n_3334), .B2 (n_3332));
AOI22_X1 i_2852 (.ZN (n_3053), .A1 (n_3488), .A2 (n_3331), .B1 (n_3329), .B2 (n_3325));
OAI21_X1 i_2851 (.ZN (n_3039), .A (n_3319), .B1 (n_3324), .B2 (n_3317));
AOI22_X1 i_2850 (.ZN (n_3032), .A1 (n_3466), .A2 (n_3316), .B1 (n_3314), .B2 (n_3312));
OAI21_X1 i_2849 (.ZN (n_3018), .A (n_3301), .B1 (n_3311), .B2 (n_3297));
OAI21_X1 i_2848 (.ZN (n_3011), .A (n_3282), .B1 (n_3292), .B2 (n_3277));
AOI21_X1 i_2847 (.ZN (n_3180), .A (n_3078), .B1 (n_3077), .B2 (n_3211));
INV_X1 i_2846 (.ZN (n_3081), .A (n_3180));
AOI21_X1 i_2845 (.ZN (n_3179), .A (n_3073), .B1 (n_3072), .B2 (n_3267));
INV_X1 i_2844 (.ZN (n_3076), .A (n_3179));
AOI21_X1 i_2843 (.ZN (n_3176), .A (n_3258), .B1 (inputB[0]), .B2 (inputA[29]));
INV_X1 i_2842 (.ZN (n_3175), .A (n_3176));
NAND3_X1 i_2841 (.ZN (n_3174), .A1 (inputB[0]), .A2 (inputA[29]), .A3 (n_3258));
NAND2_X1 i_2840 (.ZN (n_3173), .A1 (n_3175), .A2 (n_3174));
NAND2_X1 i_2839 (.ZN (n_3172), .A1 (inputB[2]), .A2 (inputA[27]));
XOR2_X1 i_2838 (.Z (n_3219), .A (n_3173), .B (n_3172));
AOI22_X1 i_2837 (.ZN (n_3171), .A1 (inputB[3]), .A2 (inputA[26]), .B1 (inputB[4]), .B2 (inputA[25]));
INV_X1 i_2836 (.ZN (n_3169), .A (n_3171));
NAND4_X1 i_2835 (.ZN (n_3168), .A1 (inputB[3]), .A2 (inputA[26]), .A3 (inputB[4]), .A4 (inputA[25]));
NAND2_X1 i_2834 (.ZN (n_3167), .A1 (n_3169), .A2 (n_3168));
NAND2_X1 i_2833 (.ZN (n_3166), .A1 (inputB[5]), .A2 (inputA[24]));
XOR2_X1 i_2832 (.Z (n_3212), .A (n_3167), .B (n_3166));
NAND2_X1 i_2831 (.ZN (n_3165), .A1 (inputB[10]), .A2 (inputA[19]));
INV_X1 i_2830 (.ZN (n_3163), .A (n_3165));
NAND2_X1 i_2829 (.ZN (n_3162), .A1 (n_3221), .A2 (n_3163));
NAND2_X1 i_2828 (.ZN (n_3161), .A1 (n_3222), .A2 (n_3165));
AND2_X1 i_2827 (.ZN (n_3160), .A1 (n_3162), .A2 (n_3161));
AND2_X1 i_2826 (.ZN (n_3159), .A1 (inputB[11]), .A2 (inputA[18]));
XOR2_X1 i_2825 (.Z (n_3198), .A (n_3160), .B (n_3159));
AOI21_X1 i_2824 (.ZN (n_3158), .A (n_3322), .B1 (inputB[13]), .B2 (inputA[16]));
INV_X1 i_2823 (.ZN (n_3155), .A (n_3158));
NAND3_X1 i_2822 (.ZN (n_3154), .A1 (inputB[13]), .A2 (inputA[16]), .A3 (n_3322));
NAND2_X1 i_2821 (.ZN (n_3150), .A1 (n_3155), .A2 (n_3154));
NAND2_X1 i_2820 (.ZN (n_3145), .A1 (inputB[14]), .A2 (inputA[15]));
XOR2_X1 i_2819 (.Z (n_3191), .A (n_3150), .B (n_3145));
NAND2_X1 i_2818 (.ZN (n_3144), .A1 (inputB[19]), .A2 (inputA[10]));
INV_X1 i_2817 (.ZN (n_3141), .A (n_3144));
NAND2_X1 i_2816 (.ZN (n_3140), .A1 (n_3196), .A2 (n_3141));
NAND2_X1 i_2815 (.ZN (n_3135), .A1 (n_3197), .A2 (n_3144));
AND2_X1 i_2814 (.ZN (n_3134), .A1 (n_3140), .A2 (n_3135));
AND2_X1 i_2813 (.ZN (n_3130), .A1 (inputB[20]), .A2 (inputA[9]));
XOR2_X1 i_2812 (.Z (n_3177), .A (n_3134), .B (n_3130));
AOI21_X1 i_2811 (.ZN (n_3125), .A (n_3302), .B1 (inputB[22]), .B2 (inputA[7]));
INV_X1 i_2810 (.ZN (n_3124), .A (n_3125));
NAND3_X1 i_2809 (.ZN (n_3120), .A1 (inputB[22]), .A2 (inputA[7]), .A3 (n_3302));
NAND2_X1 i_2808 (.ZN (n_3115), .A1 (n_3124), .A2 (n_3120));
NAND2_X1 i_2807 (.ZN (n_3114), .A1 (inputB[23]), .A2 (inputA[6]));
XOR2_X1 i_2806 (.Z (n_3170), .A (n_3115), .B (n_3114));
AOI22_X1 i_2805 (.ZN (n_3111), .A1 (inputB[27]), .A2 (inputA[2]), .B1 (inputB[28]), .B2 (inputA[1]));
INV_X1 i_2804 (.ZN (n_3110), .A (n_3111));
NAND2_X1 i_2803 (.ZN (n_3106), .A1 (inputB[28]), .A2 (inputA[2]));
INV_X1 i_2802 (.ZN (n_3105), .A (n_3106));
NAND2_X1 i_2801 (.ZN (n_3100), .A1 (n_3237), .A2 (n_3105));
NAND2_X1 i_2800 (.ZN (n_3099), .A1 (n_3110), .A2 (n_3100));
NAND2_X1 i_2799 (.ZN (n_3095), .A1 (inputB[29]), .A2 (inputA[0]));
XOR2_X1 i_2798 (.Z (n_3156), .A (n_3099), .B (n_3095));
AOI21_X1 i_2797 (.ZN (n_3091), .A (n_3083), .B1 (n_3082), .B2 (n_3271));
INV_X1 i_2796 (.ZN (n_3086), .A (n_3091));
AOI21_X1 i_2795 (.ZN (n_3090), .A (n_3200), .B1 (n_3195), .B2 (n_3192));
XOR2_X1 i_2794 (.Z (n_3231), .A (n_3229), .B (n_3090));
AOI21_X1 i_2793 (.ZN (n_3085), .A (n_3217), .B1 (n_3220), .B2 (n_3215));
XOR2_X1 i_2791 (.Z (n_3226), .A (n_3224), .B (n_3085));
AOI21_X1 i_2790 (.ZN (n_3080), .A (n_3098), .B1 (n_3097), .B2 (n_3190));
INV_X1 i_2789 (.ZN (n_3101), .A (n_3080));
AOI21_X1 i_2787 (.ZN (n_3079), .A (n_3093), .B1 (n_3092), .B2 (n_3214));
INV_X1 i_2786 (.ZN (n_3096), .A (n_3079));
AOI22_X1 i_2785 (.ZN (n_3075), .A1 (n_3403), .A2 (n_3258), .B1 (n_3252), .B2 (n_3247));
INV_X1 i_2783 (.ZN (n_3071), .A (n_3075));
XNOR2_X1 i_2782 (.ZN (n_3241), .A (n_3239), .B (n_3075));
AOI21_X1 i_2781 (.ZN (n_3070), .A (n_3113), .B1 (n_3112), .B2 (n_3203));
INV_X1 i_2779 (.ZN (n_3116), .A (n_3070));
AND2_X1 i_2778 (.ZN (n_3069), .A1 (inputB[25]), .A2 (inputA[5]));
NAND2_X1 i_2777 (.ZN (n_3068), .A1 (n_3293), .A2 (n_3069));
AOI22_X1 i_2775 (.ZN (n_3067), .A1 (inputB[24]), .A2 (inputA[5]), .B1 (inputB[25]), .B2 (inputA[4]));
INV_X1 i_2774 (.ZN (n_3066), .A (n_3067));
NAND2_X1 i_2773 (.ZN (n_3065), .A1 (n_3068), .A2 (n_3066));
NAND2_X1 i_2771 (.ZN (n_3064), .A1 (inputB[26]), .A2 (inputA[3]));
XOR2_X1 i_2770 (.Z (n_3063), .A (n_3065), .B (n_3064));
XOR2_X1 i_2769 (.Z (n_3256), .A (n_3254), .B (n_3063));
AND2_X1 i_2767 (.ZN (n_3062), .A1 (inputB[16]), .A2 (inputA[14]));
NAND2_X1 i_2766 (.ZN (n_3061), .A1 (n_3315), .A2 (n_3062));
AOI22_X1 i_2765 (.ZN (n_3058), .A1 (inputB[15]), .A2 (inputA[14]), .B1 (inputB[16]), .B2 (inputA[13]));
INV_X1 i_2763 (.ZN (n_3057), .A (n_3058));
NAND2_X1 i_2762 (.ZN (n_3056), .A1 (n_3061), .A2 (n_3057));
NAND2_X1 i_2761 (.ZN (n_3055), .A1 (inputB[17]), .A2 (inputA[12]));
XOR2_X1 i_2759 (.Z (n_3054), .A (n_3056), .B (n_3055));
XOR2_X1 i_2758 (.Z (n_3251), .A (n_3249), .B (n_3054));
AOI22_X1 i_2757 (.ZN (n_3051), .A1 (n_3364), .A2 (n_3238), .B1 (n_3236), .B2 (n_3227));
XOR2_X1 i_2755 (.Z (n_3050), .A (n_3234), .B (n_3051));
XOR2_X1 i_2754 (.Z (n_3261), .A (n_3259), .B (n_3050));
AOI21_X1 i_2753 (.ZN (n_3049), .A (n_3118), .B1 (n_3117), .B2 (n_3207));
INV_X1 i_2751 (.ZN (n_3121), .A (n_3049));
AOI21_X1 i_2750 (.ZN (n_3048), .A (n_3103), .B1 (n_3102), .B2 (n_3223));
INV_X1 i_2749 (.ZN (n_3047), .A (n_3048));
XNOR2_X1 i_2747 (.ZN (n_3266), .A (n_3264), .B (n_3048));
AOI21_X1 i_2746 (.ZN (n_3046), .A (n_3123), .B1 (n_3122), .B2 (n_3189));
INV_X1 i_2745 (.ZN (n_3126), .A (n_3046));
AOI21_X1 i_2743 (.ZN (n_3045), .A (n_3128), .B1 (n_3127), .B2 (n_3202));
INV_X1 i_2742 (.ZN (n_3131), .A (n_3045));
AOI21_X1 i_2741 (.ZN (n_3044), .A (n_3133), .B1 (n_3132), .B2 (n_3183));
INV_X1 i_2739 (.ZN (n_3136), .A (n_3044));
AOI21_X1 i_2738 (.ZN (n_3043), .A (n_3088), .B1 (n_3087), .B2 (n_3246));
INV_X1 i_2737 (.ZN (n_3042), .A (n_3043));
XNOR2_X1 i_2735 (.ZN (n_3041), .A (n_3269), .B (n_3043));
XOR2_X1 i_2734 (.Z (n_3286), .A (n_3284), .B (n_3041));
AOI21_X1 i_2733 (.ZN (n_3040), .A (n_3108), .B1 (n_3107), .B2 (n_3210));
INV_X1 i_2731 (.ZN (n_3037), .A (n_3040));
XNOR2_X1 i_2730 (.ZN (n_3036), .A (n_3274), .B (n_3040));
XOR2_X1 i_2729 (.Z (n_3291), .A (n_3289), .B (n_3036));
AOI21_X1 i_2728 (.ZN (n_3035), .A (n_3143), .B1 (n_3142), .B2 (n_3182));
INV_X1 i_2727 (.ZN (n_3146), .A (n_3035));
AND2_X1 i_2726 (.ZN (n_3034), .A1 (inputB[7]), .A2 (inputA[23]));
NAND2_X1 i_2725 (.ZN (n_3033), .A1 (n_3330), .A2 (n_3034));
AOI22_X1 i_2724 (.ZN (n_3030), .A1 (inputB[6]), .A2 (inputA[23]), .B1 (inputB[7]), .B2 (inputA[22]));
INV_X1 i_2723 (.ZN (n_3029), .A (n_3030));
NAND2_X1 i_2722 (.ZN (n_3028), .A1 (n_3033), .A2 (n_3029));
NAND2_X1 i_2721 (.ZN (n_3027), .A1 (inputB[8]), .A2 (inputA[21]));
XOR2_X1 i_2720 (.Z (n_3026), .A (n_3028), .B (n_3027));
XOR2_X1 i_2719 (.Z (n_3025), .A (n_3244), .B (n_3026));
XOR2_X1 i_2718 (.Z (n_3024), .A (n_3279), .B (n_3025));
XOR2_X1 i_2717 (.Z (n_3296), .A (n_3294), .B (n_3024));
AOI21_X1 i_2716 (.ZN (n_3023), .A (n_3148), .B1 (n_3147), .B2 (n_3181));
INV_X1 i_2715 (.ZN (n_3151), .A (n_3023));
AOI21_X1 i_2714 (.ZN (n_3022), .A (n_3138), .B1 (n_3137), .B2 (n_3188));
INV_X1 i_2713 (.ZN (n_3021), .A (n_3022));
XNOR2_X1 i_2712 (.ZN (n_3020), .A (n_3299), .B (n_3022));
XOR2_X1 i_2711 (.Z (n_3306), .A (n_3304), .B (n_3020));
OAI21_X1 i_2710 (.ZN (n_3206), .A (n_3033), .B1 (n_3030), .B2 (n_3027));
NAND2_X1 i_2709 (.ZN (n_3019), .A1 (n_3161), .A2 (n_3159));
NAND2_X1 i_2708 (.ZN (n_3199), .A1 (n_3162), .A2 (n_3019));
OAI21_X1 i_2707 (.ZN (n_3185), .A (n_3061), .B1 (n_3058), .B2 (n_3055));
NAND2_X1 i_2706 (.ZN (n_3016), .A1 (n_3135), .A2 (n_3130));
NAND2_X1 i_2705 (.ZN (n_3178), .A1 (n_3140), .A2 (n_3016));
OAI21_X1 i_2704 (.ZN (n_3164), .A (n_3068), .B1 (n_3067), .B2 (n_3064));
OAI21_X1 i_2703 (.ZN (n_3157), .A (n_3100), .B1 (n_3111), .B2 (n_3095));
AOI21_X1 i_2702 (.ZN (n_3015), .A (n_3230), .B1 (n_3229), .B2 (n_3090));
INV_X1 i_2701 (.ZN (n_3233), .A (n_3015));
AOI21_X1 i_2700 (.ZN (n_3014), .A (n_3225), .B1 (n_3224), .B2 (n_3085));
INV_X1 i_2699 (.ZN (n_3228), .A (n_3014));
AND2_X1 i_2698 (.ZN (n_3013), .A1 (inputB[5]), .A2 (inputA[25]));
AOI21_X1 i_2697 (.ZN (n_3012), .A (n_3013), .B1 (inputB[4]), .B2 (inputA[26]));
INV_X1 i_2696 (.ZN (n_3009), .A (n_3012));
NAND3_X1 i_2695 (.ZN (n_3008), .A1 (inputB[4]), .A2 (inputA[26]), .A3 (n_3013));
NAND2_X1 i_2694 (.ZN (n_3007), .A1 (n_3009), .A2 (n_3008));
NAND2_X1 i_2693 (.ZN (n_3006), .A1 (inputB[6]), .A2 (inputA[24]));
XOR2_X1 i_2692 (.Z (n_3369), .A (n_3007), .B (n_3006));
AOI21_X1 i_2691 (.ZN (n_3005), .A (n_3034), .B1 (inputB[8]), .B2 (inputA[22]));
INV_X1 i_2690 (.ZN (n_3004), .A (n_3005));
NAND3_X1 i_2689 (.ZN (n_3003), .A1 (inputB[8]), .A2 (inputA[22]), .A3 (n_3034));
NAND2_X1 i_2688 (.ZN (n_3002), .A1 (n_3004), .A2 (n_3003));
NAND2_X1 i_2687 (.ZN (n_3001), .A1 (inputB[9]), .A2 (inputA[21]));
XOR2_X1 i_2686 (.Z (n_3362), .A (n_3002), .B (n_3001));
AND2_X1 i_2685 (.ZN (n_2997), .A1 (inputB[14]), .A2 (inputA[16]));
NAND3_X1 i_2684 (.ZN (n_2992), .A1 (inputB[13]), .A2 (inputA[17]), .A3 (n_2997));
INV_X1 i_2683 (.ZN (n_2991), .A (n_2992));
AOI21_X1 i_2682 (.ZN (n_2987), .A (n_2997), .B1 (inputB[13]), .B2 (inputA[17]));
NOR2_X1 i_2681 (.ZN (n_2982), .A1 (n_2991), .A2 (n_2987));
NAND2_X1 i_2680 (.ZN (n_2981), .A1 (inputB[15]), .A2 (inputA[15]));
XNOR2_X1 i_2679 (.ZN (n_3348), .A (n_2982), .B (n_2981));
AOI21_X1 i_2678 (.ZN (n_2978), .A (n_3062), .B1 (inputB[17]), .B2 (inputA[13]));
INV_X1 i_2677 (.ZN (n_2977), .A (n_2978));
NAND3_X1 i_2676 (.ZN (n_2972), .A1 (inputB[17]), .A2 (inputA[13]), .A3 (n_3062));
NAND2_X1 i_2675 (.ZN (n_2967), .A1 (n_2977), .A2 (n_2972));
NAND2_X1 i_2674 (.ZN (n_2963), .A1 (inputB[18]), .A2 (inputA[12]));
XOR2_X1 i_2673 (.Z (n_3341), .A (n_2967), .B (n_2963));
AND2_X1 i_2672 (.ZN (n_2962), .A1 (inputB[23]), .A2 (inputA[7]));
AOI21_X1 i_2671 (.ZN (n_2957), .A (n_2962), .B1 (inputB[22]), .B2 (inputA[8]));
INV_X1 i_2670 (.ZN (n_2952), .A (n_2957));
NAND3_X1 i_2669 (.ZN (n_2951), .A1 (inputB[22]), .A2 (inputA[8]), .A3 (n_2962));
NAND2_X1 i_2668 (.ZN (n_2948), .A1 (n_2952), .A2 (n_2951));
NAND2_X1 i_2667 (.ZN (n_2947), .A1 (inputB[24]), .A2 (inputA[6]));
XOR2_X1 i_2666 (.Z (n_3327), .A (n_2948), .B (n_2947));
AOI21_X1 i_2665 (.ZN (n_2942), .A (n_3069), .B1 (inputB[26]), .B2 (inputA[4]));
INV_X1 i_2664 (.ZN (n_2937), .A (n_2942));
NAND3_X1 i_2663 (.ZN (n_2936), .A1 (inputB[26]), .A2 (inputA[4]), .A3 (n_3069));
NAND2_X1 i_2662 (.ZN (n_2933), .A1 (n_2937), .A2 (n_2936));
NAND2_X1 i_2661 (.ZN (n_2932), .A1 (inputB[27]), .A2 (inputA[3]));
XOR2_X1 i_2659 (.Z (n_3320), .A (n_2933), .B (n_2932));
AOI21_X1 i_2658 (.ZN (n_2927), .A (n_3240), .B1 (n_3239), .B2 (n_3071));
INV_X1 i_2657 (.ZN (n_3243), .A (n_2927));
AOI21_X1 i_2655 (.ZN (n_2926), .A (n_3235), .B1 (n_3234), .B2 (n_3051));
INV_X1 i_2654 (.ZN (n_2923), .A (n_2926));
XNOR2_X1 i_2653 (.ZN (n_3401), .A (n_3399), .B (n_2926));
OAI21_X1 i_2651 (.ZN (n_2922), .A (n_3154), .B1 (n_3158), .B2 (n_3145));
XOR2_X1 i_2650 (.Z (n_3391), .A (n_3389), .B (n_2922));
OAI21_X1 i_2649 (.ZN (n_2921), .A (n_3174), .B1 (n_3176), .B2 (n_3172));
OAI21_X1 i_2647 (.ZN (n_2920), .A (n_3168), .B1 (n_3171), .B2 (n_3166));
NAND2_X1 i_2646 (.ZN (n_2917), .A1 (n_2921), .A2 (n_2920));
NOR2_X1 i_2645 (.ZN (n_2916), .A1 (n_2921), .A2 (n_2920));
AOI21_X1 i_2643 (.ZN (n_2915), .A (n_2916), .B1 (n_2921), .B2 (n_2920));
NAND2_X1 i_2642 (.ZN (n_2914), .A1 (inputB[0]), .A2 (inputA[30]));
XNOR2_X1 i_2641 (.ZN (n_3383), .A (n_2915), .B (n_2914));
AOI21_X1 i_2639 (.ZN (n_2913), .A (n_3250), .B1 (n_3249), .B2 (n_3054));
INV_X1 i_2638 (.ZN (n_3253), .A (n_2913));
AOI21_X1 i_2637 (.ZN (n_2912), .A (n_3245), .B1 (n_3244), .B2 (n_3026));
INV_X1 i_2635 (.ZN (n_3248), .A (n_2912));
AOI21_X1 i_2634 (.ZN (n_2910), .A (n_3270), .B1 (n_3269), .B2 (n_3042));
INV_X1 i_2633 (.ZN (n_3273), .A (n_2910));
AOI21_X1 i_2631 (.ZN (n_2909), .A (n_3265), .B1 (n_3264), .B2 (n_3047));
INV_X1 i_2630 (.ZN (n_3268), .A (n_2909));
NAND2_X1 i_2629 (.ZN (n_2908), .A1 (inputB[29]), .A2 (inputA[1]));
INV_X1 i_2627 (.ZN (n_2907), .A (n_2908));
NAND2_X1 i_2626 (.ZN (n_2906), .A1 (n_3105), .A2 (n_2907));
OAI21_X1 i_2625 (.ZN (n_2903), .A (n_2906), .B1 (n_3105), .B2 (n_2907));
NAND2_X1 i_2623 (.ZN (n_2902), .A1 (inputB[30]), .A2 (inputA[0]));
XOR2_X1 i_2622 (.Z (n_2901), .A (n_2903), .B (n_2902));
XOR2_X1 i_2621 (.Z (n_3421), .A (n_3419), .B (n_2901));
NAND2_X1 i_2619 (.ZN (n_2900), .A1 (inputB[20]), .A2 (inputA[11]));
INV_X1 i_2618 (.ZN (n_2899), .A (n_2900));
NAND2_X1 i_2617 (.ZN (n_2897), .A1 (n_3141), .A2 (n_2899));
AOI22_X1 i_2615 (.ZN (n_2896), .A1 (inputB[19]), .A2 (inputA[11]), .B1 (inputB[20]), .B2 (inputA[10]));
INV_X1 i_2614 (.ZN (n_2895), .A (n_2896));
NAND2_X1 i_2613 (.ZN (n_2894), .A1 (n_2897), .A2 (n_2895));
NAND2_X1 i_2611 (.ZN (n_2893), .A1 (inputB[21]), .A2 (inputA[9]));
XOR2_X1 i_2610 (.Z (n_2892), .A (n_2894), .B (n_2893));
XOR2_X1 i_2609 (.Z (n_3416), .A (n_3414), .B (n_2892));
AOI21_X1 i_2607 (.ZN (n_2891), .A (n_3275), .B1 (n_3274), .B2 (n_3037));
INV_X1 i_2606 (.ZN (n_3278), .A (n_2891));
NAND2_X1 i_2605 (.ZN (n_2889), .A1 (inputB[2]), .A2 (inputA[29]));
NAND3_X1 i_2603 (.ZN (n_2888), .A1 (inputB[2]), .A2 (inputA[29]), .A3 (n_3258));
AOI22_X1 i_2602 (.ZN (n_2887), .A1 (inputB[1]), .A2 (inputA[29]), .B1 (inputB[2]), .B2 (inputA[28]));
INV_X1 i_2601 (.ZN (n_2886), .A (n_2887));
NAND2_X1 i_2599 (.ZN (n_2885), .A1 (n_2888), .A2 (n_2886));
NAND2_X1 i_2598 (.ZN (n_2882), .A1 (inputB[3]), .A2 (inputA[27]));
XOR2_X1 i_2597 (.Z (n_2881), .A (n_2885), .B (n_2882));
XOR2_X1 i_2596 (.Z (n_2880), .A (n_3404), .B (n_2881));
XOR2_X1 i_2595 (.Z (n_3436), .A (n_3434), .B (n_2880));
OAI21_X1 i_2594 (.ZN (n_2879), .A (n_3120), .B1 (n_3125), .B2 (n_3114));
XOR2_X1 i_2593 (.Z (n_2878), .A (n_3394), .B (n_2879));
XOR2_X1 i_2592 (.Z (n_3426), .A (n_3424), .B (n_2878));
AOI21_X1 i_2591 (.ZN (n_2876), .A (n_3280), .B1 (n_3279), .B2 (n_3025));
INV_X1 i_2590 (.ZN (n_3283), .A (n_2876));
AOI21_X1 i_2589 (.ZN (n_2875), .A (n_3285), .B1 (n_3284), .B2 (n_3041));
INV_X1 i_2588 (.ZN (n_3288), .A (n_2875));
AOI22_X1 i_2587 (.ZN (n_2874), .A1 (inputB[10]), .A2 (inputA[20]), .B1 (inputB[11]), .B2 (inputA[19]));
INV_X1 i_2586 (.ZN (n_2873), .A (n_2874));
NAND2_X1 i_2585 (.ZN (n_2872), .A1 (inputB[11]), .A2 (inputA[20]));
INV_X1 i_2584 (.ZN (n_2871), .A (n_2872));
NAND2_X1 i_2583 (.ZN (n_2870), .A1 (n_3163), .A2 (n_2871));
NAND2_X1 i_2582 (.ZN (n_2868), .A1 (n_2873), .A2 (n_2870));
NAND2_X1 i_2581 (.ZN (n_2867), .A1 (inputB[12]), .A2 (inputA[18]));
XOR2_X1 i_2580 (.Z (n_2866), .A (n_2868), .B (n_2867));
XOR2_X1 i_2579 (.Z (n_2865), .A (n_3409), .B (n_2866));
XOR2_X1 i_2578 (.Z (n_3446), .A (n_3444), .B (n_2865));
AOI21_X1 i_2577 (.ZN (n_2864), .A (n_3260), .B1 (n_3259), .B2 (n_3050));
INV_X1 i_2576 (.ZN (n_2861), .A (n_2864));
XNOR2_X1 i_2575 (.ZN (n_2860), .A (n_3439), .B (n_2864));
XOR2_X1 i_2574 (.Z (n_3456), .A (n_3454), .B (n_2860));
AOI21_X1 i_2573 (.ZN (n_2859), .A (n_3255), .B1 (n_3254), .B2 (n_3063));
INV_X1 i_2572 (.ZN (n_2858), .A (n_2859));
XNOR2_X1 i_2571 (.ZN (n_2857), .A (n_3429), .B (n_2859));
XOR2_X1 i_2570 (.Z (n_3451), .A (n_3449), .B (n_2857));
AOI21_X1 i_2569 (.ZN (n_2855), .A (n_3300), .B1 (n_3299), .B2 (n_3021));
INV_X1 i_2568 (.ZN (n_3303), .A (n_2855));
AOI21_X1 i_2567 (.ZN (n_2854), .A (n_3290), .B1 (n_3289), .B2 (n_3036));
INV_X1 i_2566 (.ZN (n_2853), .A (n_2854));
XNOR2_X1 i_2565 (.ZN (n_3461), .A (n_3459), .B (n_2854));
AOI21_X1 i_2564 (.ZN (n_2849), .A (n_3305), .B1 (n_3304), .B2 (n_3020));
INV_X1 i_2563 (.ZN (n_3308), .A (n_2849));
AOI21_X1 i_2562 (.ZN (n_2844), .A (n_3295), .B1 (n_3294), .B2 (n_3024));
INV_X1 i_2561 (.ZN (n_2843), .A (n_2844));
XNOR2_X1 i_2560 (.ZN (n_2839), .A (n_3464), .B (n_2844));
XOR2_X1 i_2559 (.Z (n_3471), .A (n_3469), .B (n_2839));
OAI21_X1 i_2558 (.ZN (n_3370), .A (n_3008), .B1 (n_3012), .B2 (n_3006));
OAI21_X1 i_2557 (.ZN (n_3363), .A (n_3003), .B1 (n_3005), .B2 (n_3001));
OAI21_X1 i_2556 (.ZN (n_3349), .A (n_2992), .B1 (n_2987), .B2 (n_2981));
OAI21_X1 i_2555 (.ZN (n_3342), .A (n_2972), .B1 (n_2978), .B2 (n_2963));
OAI21_X1 i_2554 (.ZN (n_3328), .A (n_2951), .B1 (n_2957), .B2 (n_2947));
OAI21_X1 i_2553 (.ZN (n_3321), .A (n_2936), .B1 (n_2942), .B2 (n_2932));
AOI21_X1 i_2552 (.ZN (n_2835), .A (n_3395), .B1 (n_3394), .B2 (n_2879));
INV_X1 i_2551 (.ZN (n_3398), .A (n_2835));
AOI21_X1 i_2550 (.ZN (n_2834), .A (n_3390), .B1 (n_3389), .B2 (n_2922));
INV_X1 i_2549 (.ZN (n_3393), .A (n_2834));
OAI211_X1 i_2548 (.ZN (n_2833), .A (inputB[0]), .B (inputA[31]), .C1 (n_5754), .C2 (n_5751));
AOI211_X1 i_2547 (.ZN (n_2830), .A (n_5754), .B (n_5751), .C1 (inputB[0]), .C2 (inputA[31]));
INV_X1 i_2546 (.ZN (n_2829), .A (n_2830));
NAND2_X1 i_2545 (.ZN (n_2825), .A1 (n_2833), .A2 (n_2829));
OAI21_X1 i_2544 (.ZN (n_2824), .A (n_2888), .B1 (n_2887), .B2 (n_2882));
XNOR2_X1 i_2543 (.ZN (n_3549), .A (n_2825), .B (n_2824));
NAND2_X1 i_2542 (.ZN (n_2819), .A1 (inputB[3]), .A2 (inputA[28]));
OR2_X1 i_2541 (.ZN (n_2814), .A1 (n_2889), .A2 (n_2819));
NAND2_X1 i_2540 (.ZN (n_2813), .A1 (n_2889), .A2 (n_2819));
AND2_X1 i_2539 (.ZN (n_2809), .A1 (n_2814), .A2 (n_2813));
NAND2_X1 i_2538 (.ZN (n_2804), .A1 (inputB[4]), .A2 (inputA[27]));
XNOR2_X1 i_2537 (.ZN (n_3542), .A (n_2809), .B (n_2804));
AND2_X1 i_2535 (.ZN (n_2800), .A1 (inputB[9]), .A2 (inputA[22]));
AOI21_X1 i_2534 (.ZN (n_2799), .A (n_2800), .B1 (inputB[8]), .B2 (inputA[23]));
INV_X1 i_2533 (.ZN (n_2798), .A (n_2799));
NAND3_X1 i_2531 (.ZN (n_2794), .A1 (inputB[8]), .A2 (inputA[23]), .A3 (n_2800));
NAND2_X1 i_2530 (.ZN (n_2789), .A1 (n_2798), .A2 (n_2794));
NAND2_X1 i_2529 (.ZN (n_2784), .A1 (inputB[10]), .A2 (inputA[21]));
XOR2_X1 i_2527 (.Z (n_3528), .A (n_2789), .B (n_2784));
NAND2_X1 i_2526 (.ZN (n_2780), .A1 (inputB[12]), .A2 (inputA[19]));
INV_X1 i_2525 (.ZN (n_2779), .A (n_2780));
NAND2_X1 i_2523 (.ZN (n_2778), .A1 (n_2871), .A2 (n_2779));
OAI21_X1 i_2522 (.ZN (n_2775), .A (n_2778), .B1 (n_2871), .B2 (n_2779));
NAND2_X1 i_2521 (.ZN (n_2774), .A1 (inputB[13]), .A2 (inputA[18]));
XOR2_X1 i_2519 (.Z (n_3521), .A (n_2775), .B (n_2774));
AND2_X1 i_2518 (.ZN (n_2773), .A1 (inputB[18]), .A2 (inputA[13]));
AOI21_X1 i_2517 (.ZN (n_2772), .A (n_2773), .B1 (inputB[17]), .B2 (inputA[14]));
INV_X1 i_2515 (.ZN (n_2771), .A (n_2772));
NAND3_X1 i_2514 (.ZN (n_2770), .A1 (inputB[17]), .A2 (inputA[14]), .A3 (n_2773));
NAND2_X1 i_2513 (.ZN (n_2769), .A1 (n_2771), .A2 (n_2770));
NAND2_X1 i_2511 (.ZN (n_2768), .A1 (inputB[19]), .A2 (inputA[12]));
XOR2_X1 i_2510 (.Z (n_3507), .A (n_2769), .B (n_2768));
NAND2_X1 i_2509 (.ZN (n_2767), .A1 (inputB[21]), .A2 (inputA[10]));
INV_X1 i_2507 (.ZN (n_2766), .A (n_2767));
NAND2_X1 i_2506 (.ZN (n_2765), .A1 (n_2899), .A2 (n_2766));
NAND2_X1 i_2505 (.ZN (n_2763), .A1 (n_2900), .A2 (n_2767));
AND2_X1 i_2503 (.ZN (n_2762), .A1 (n_2765), .A2 (n_2763));
AND2_X1 i_2502 (.ZN (n_2761), .A1 (inputB[22]), .A2 (inputA[9]));
XOR2_X1 i_2501 (.Z (n_3500), .A (n_2762), .B (n_2761));
AND2_X1 i_2499 (.ZN (n_2760), .A1 (inputB[27]), .A2 (inputA[4]));
AOI21_X1 i_2498 (.ZN (n_2759), .A (n_2760), .B1 (inputB[26]), .B2 (inputA[5]));
INV_X1 i_2497 (.ZN (n_2756), .A (n_2759));
NAND3_X1 i_2495 (.ZN (n_2755), .A1 (inputB[26]), .A2 (inputA[5]), .A3 (n_2760));
NAND2_X1 i_2494 (.ZN (n_2754), .A1 (n_2756), .A2 (n_2755));
NAND2_X1 i_2493 (.ZN (n_2753), .A1 (inputB[28]), .A2 (inputA[3]));
XOR2_X1 i_2491 (.Z (n_3486), .A (n_2754), .B (n_2753));
AOI22_X1 i_2490 (.ZN (n_2752), .A1 (inputB[29]), .A2 (inputA[2]), .B1 (inputB[30]), .B2 (inputA[1]));
INV_X1 i_2489 (.ZN (n_2750), .A (n_2752));
NAND2_X1 i_2487 (.ZN (n_2749), .A1 (inputB[30]), .A2 (inputA[2]));
OR2_X1 i_2486 (.ZN (n_2748), .A1 (n_2908), .A2 (n_2749));
NAND2_X1 i_2485 (.ZN (n_2747), .A1 (n_2750), .A2 (n_2748));
NAND2_X1 i_2483 (.ZN (n_2746), .A1 (inputB[31]), .A2 (inputA[0]));
INV_X1 i_2482 (.ZN (n_2745), .A (n_2746));
XNOR2_X1 i_2481 (.ZN (n_3477), .A (n_2747), .B (n_2746));
AOI22_X1 i_2479 (.ZN (n_2744), .A1 (n_3106), .A2 (n_2908), .B1 (n_2906), .B2 (n_2902));
XOR2_X1 i_2478 (.Z (n_3567), .A (n_3565), .B (n_2744));
AOI21_X1 i_2477 (.ZN (n_2742), .A (n_2896), .B1 (n_2897), .B2 (n_2893));
XOR2_X1 i_2476 (.Z (n_3562), .A (n_3560), .B (n_2742));
AOI21_X1 i_2475 (.ZN (n_2741), .A (n_3420), .B1 (n_3419), .B2 (n_2901));
INV_X1 i_2474 (.ZN (n_3423), .A (n_2741));
AOI21_X1 i_2473 (.ZN (n_2740), .A (n_3415), .B1 (n_3414), .B2 (n_2892));
INV_X1 i_2472 (.ZN (n_3418), .A (n_2740));
AOI21_X1 i_2471 (.ZN (n_2739), .A (n_3405), .B1 (n_3404), .B2 (n_2881));
INV_X1 i_2470 (.ZN (n_3408), .A (n_2739));
OAI21_X1 i_2469 (.ZN (n_2738), .A (n_2917), .B1 (n_2916), .B2 (n_2914));
XOR2_X1 i_2468 (.Z (n_3572), .A (n_3570), .B (n_2738));
AOI21_X1 i_2467 (.ZN (n_2735), .A (n_3425), .B1 (n_3424), .B2 (n_2878));
INV_X1 i_2466 (.ZN (n_3428), .A (n_2735));
AOI21_X1 i_2465 (.ZN (n_2734), .A (n_3400), .B1 (n_3399), .B2 (n_2923));
INV_X1 i_2464 (.ZN (n_2733), .A (n_2734));
XNOR2_X1 i_2463 (.ZN (n_3592), .A (n_3590), .B (n_2734));
NAND3_X1 i_2462 (.ZN (n_2732), .A1 (inputB[15]), .A2 (inputA[17]), .A3 (n_2997));
AOI22_X1 i_2461 (.ZN (n_2731), .A1 (inputB[14]), .A2 (inputA[17]), .B1 (inputB[15]), .B2 (inputA[16]));
INV_X1 i_2460 (.ZN (n_2729), .A (n_2731));
NAND2_X1 i_2459 (.ZN (n_2728), .A1 (n_2732), .A2 (n_2729));
NAND2_X1 i_2458 (.ZN (n_2727), .A1 (inputB[16]), .A2 (inputA[15]));
XOR2_X1 i_2457 (.Z (n_2726), .A (n_2728), .B (n_2727));
XOR2_X1 i_2456 (.Z (n_3582), .A (n_3580), .B (n_2726));
NAND3_X1 i_2455 (.ZN (n_2725), .A1 (inputB[6]), .A2 (inputA[26]), .A3 (n_3013));
AOI22_X1 i_2454 (.ZN (n_2724), .A1 (inputB[5]), .A2 (inputA[26]), .B1 (inputB[6]), .B2 (inputA[25]));
INV_X1 i_2453 (.ZN (n_2723), .A (n_2724));
NAND2_X1 i_2452 (.ZN (n_2721), .A1 (n_2725), .A2 (n_2723));
NAND2_X1 i_2451 (.ZN (n_2720), .A1 (inputB[7]), .A2 (inputA[24]));
XOR2_X1 i_2450 (.Z (n_2719), .A (n_2721), .B (n_2720));
XOR2_X1 i_2449 (.Z (n_3577), .A (n_3575), .B (n_2719));
AOI21_X1 i_2448 (.ZN (n_2718), .A (n_3435), .B1 (n_3434), .B2 (n_2880));
INV_X1 i_2447 (.ZN (n_3438), .A (n_2718));
AOI21_X1 i_2446 (.ZN (n_2717), .A (n_3410), .B1 (n_3409), .B2 (n_2866));
INV_X1 i_2445 (.ZN (n_2714), .A (n_2717));
XNOR2_X1 i_2444 (.ZN (n_3602), .A (n_3600), .B (n_2717));
AOI21_X1 i_2443 (.ZN (n_2713), .A (n_3445), .B1 (n_3444), .B2 (n_2865));
INV_X1 i_2442 (.ZN (n_3448), .A (n_2713));
AOI21_X1 i_2441 (.ZN (n_2709), .A (n_3430), .B1 (n_3429), .B2 (n_2858));
INV_X1 i_2440 (.ZN (n_2704), .A (n_2709));
XNOR2_X1 i_2439 (.ZN (n_3607), .A (n_3605), .B (n_2709));
AOI21_X1 i_2438 (.ZN (n_2703), .A (n_3440), .B1 (n_3439), .B2 (n_2861));
INV_X1 i_2437 (.ZN (n_2699), .A (n_2703));
XNOR2_X1 i_2436 (.ZN (n_3617), .A (n_3615), .B (n_2703));
NAND3_X1 i_2435 (.ZN (n_2695), .A1 (inputB[24]), .A2 (inputA[8]), .A3 (n_2962));
AOI22_X1 i_2434 (.ZN (n_2694), .A1 (inputB[23]), .A2 (inputA[8]), .B1 (inputB[24]), .B2 (inputA[7]));
INV_X1 i_2433 (.ZN (n_2693), .A (n_2694));
NAND2_X1 i_2432 (.ZN (n_2689), .A1 (n_2695), .A2 (n_2693));
NAND2_X1 i_2431 (.ZN (n_2684), .A1 (inputB[25]), .A2 (inputA[6]));
XOR2_X1 i_2430 (.Z (n_2679), .A (n_2689), .B (n_2684));
XOR2_X1 i_2429 (.Z (n_2675), .A (n_3585), .B (n_2679));
XOR2_X1 i_2428 (.Z (n_3612), .A (n_3610), .B (n_2675));
OAI21_X1 i_2427 (.ZN (n_2674), .A (n_2870), .B1 (n_2874), .B2 (n_2867));
XOR2_X1 i_2426 (.Z (n_2673), .A (n_3555), .B (n_2674));
XOR2_X1 i_2425 (.Z (n_2669), .A (n_3595), .B (n_2673));
XOR2_X1 i_2424 (.Z (n_3622), .A (n_3620), .B (n_2669));
AOI21_X1 i_2423 (.ZN (n_2664), .A (n_3460), .B1 (n_3459), .B2 (n_2853));
INV_X1 i_2422 (.ZN (n_3463), .A (n_2664));
AOI21_X1 i_2421 (.ZN (n_2660), .A (n_3465), .B1 (n_3464), .B2 (n_2843));
INV_X1 i_2420 (.ZN (n_3468), .A (n_2660));
AOI21_X1 i_2419 (.ZN (n_2659), .A (n_3455), .B1 (n_3454), .B2 (n_2860));
INV_X1 i_2418 (.ZN (n_2658), .A (n_2659));
XNOR2_X1 i_2417 (.ZN (n_3632), .A (n_3630), .B (n_2659));
AOI21_X1 i_2416 (.ZN (n_2655), .A (n_3470), .B1 (n_3469), .B2 (n_2839));
INV_X1 i_2414 (.ZN (n_3473), .A (n_2655));
AOI21_X1 i_2413 (.ZN (n_2654), .A (n_3450), .B1 (n_3449), .B2 (n_2857));
INV_X1 i_2412 (.ZN (n_2650), .A (n_2654));
XNOR2_X1 i_2410 (.ZN (n_2649), .A (n_3625), .B (n_2654));
XOR2_X1 i_2409 (.Z (n_2644), .A (n_3635), .B (n_2649));
XOR2_X1 i_2408 (.Z (n_3642), .A (n_3640), .B (n_2644));
OAI21_X1 i_2406 (.ZN (n_3536), .A (n_2725), .B1 (n_2724), .B2 (n_2720));
OAI21_X1 i_2405 (.ZN (n_3529), .A (n_2794), .B1 (n_2799), .B2 (n_2784));
OAI21_X1 i_2404 (.ZN (n_3515), .A (n_2732), .B1 (n_2731), .B2 (n_2727));
OAI21_X1 i_2402 (.ZN (n_3508), .A (n_2770), .B1 (n_2772), .B2 (n_2768));
OAI21_X1 i_2401 (.ZN (n_3494), .A (n_2695), .B1 (n_2694), .B2 (n_2684));
OAI21_X1 i_2400 (.ZN (n_3487), .A (n_2755), .B1 (n_2759), .B2 (n_2753));
AOI21_X1 i_2398 (.ZN (n_2643), .A (n_3566), .B1 (n_3565), .B2 (n_2744));
INV_X1 i_2397 (.ZN (n_3569), .A (n_2643));
AOI21_X1 i_2396 (.ZN (n_2640), .A (n_3561), .B1 (n_3560), .B2 (n_2742));
INV_X1 i_2394 (.ZN (n_3564), .A (n_2640));
AOI21_X1 i_2393 (.ZN (n_2639), .A (n_2830), .B1 (n_2833), .B2 (n_2824));
INV_X1 i_2392 (.ZN (n_3550), .A (n_2639));
OAI211_X1 i_2390 (.ZN (n_2638), .A (inputB[1]), .B (inputA[31]), .C1 (n_5755), .C2 (n_5751));
OAI211_X1 i_2389 (.ZN (n_2637), .A (inputB[2]), .B (inputA[30]), .C1 (n_5754), .C2 (n_5753));
NAND2_X1 i_2388 (.ZN (n_2636), .A1 (n_2814), .A2 (n_2804));
NAND2_X1 i_2386 (.ZN (n_2633), .A1 (n_2813), .A2 (n_2636));
AOI21_X1 i_2385 (.ZN (n_2632), .A (n_2633), .B1 (n_2638), .B2 (n_2637));
NAND2_X1 i_2384 (.ZN (n_2631), .A1 (n_2637), .A2 (n_2633));
INV_X1 i_2382 (.ZN (n_2630), .A (n_2631));
AOI21_X1 i_2381 (.ZN (n_2628), .A (n_2632), .B1 (n_2638), .B2 (n_2630));
INV_X1 i_2380 (.ZN (n_3716), .A (n_2628));
AOI22_X1 i_2378 (.ZN (n_2627), .A1 (inputB[6]), .A2 (inputA[26]), .B1 (inputB[7]), .B2 (inputA[25]));
INV_X1 i_2377 (.ZN (n_2626), .A (n_2627));
NAND2_X1 i_2376 (.ZN (n_2625), .A1 (inputB[7]), .A2 (inputA[26]));
INV_X1 i_2374 (.ZN (n_2624), .A (n_2625));
NAND3_X1 i_2373 (.ZN (n_2623), .A1 (inputB[6]), .A2 (inputA[25]), .A3 (n_2624));
NAND2_X1 i_2372 (.ZN (n_2620), .A1 (n_2626), .A2 (n_2623));
NAND2_X1 i_2370 (.ZN (n_2619), .A1 (inputB[8]), .A2 (inputA[24]));
XOR2_X1 i_2369 (.Z (n_3702), .A (n_2620), .B (n_2619));
AND2_X1 i_2368 (.ZN (n_2618), .A1 (inputB[10]), .A2 (inputA[23]));
NAND2_X1 i_2366 (.ZN (n_2617), .A1 (n_2800), .A2 (n_2618));
AOI22_X1 i_2365 (.ZN (n_2616), .A1 (inputB[9]), .A2 (inputA[23]), .B1 (inputB[10]), .B2 (inputA[22]));
INV_X1 i_2364 (.ZN (n_2615), .A (n_2616));
NAND2_X1 i_2362 (.ZN (n_2613), .A1 (n_2617), .A2 (n_2615));
NAND2_X1 i_2361 (.ZN (n_2612), .A1 (inputB[11]), .A2 (inputA[21]));
XOR2_X1 i_2360 (.Z (n_3695), .A (n_2613), .B (n_2612));
NAND2_X1 i_2359 (.ZN (n_2611), .A1 (inputB[17]), .A2 (inputA[15]));
INV_X1 i_2358 (.ZN (n_2610), .A (n_2611));
AOI22_X1 i_2357 (.ZN (n_2609), .A1 (inputB[15]), .A2 (inputA[17]), .B1 (inputB[16]), .B2 (inputA[16]));
AND2_X1 i_2356 (.ZN (n_2607), .A1 (inputB[16]), .A2 (inputA[17]));
NAND3_X1 i_2355 (.ZN (n_2606), .A1 (inputB[15]), .A2 (inputA[16]), .A3 (n_2607));
INV_X1 i_2354 (.ZN (n_2605), .A (n_2606));
NOR2_X1 i_2353 (.ZN (n_2604), .A1 (n_2609), .A2 (n_2605));
XOR2_X1 i_2352 (.Z (n_3681), .A (n_2610), .B (n_2604));
NAND2_X1 i_2351 (.ZN (n_2603), .A1 (inputB[19]), .A2 (inputA[14]));
INV_X1 i_2350 (.ZN (n_2602), .A (n_2603));
NAND2_X1 i_2349 (.ZN (n_2599), .A1 (n_2773), .A2 (n_2602));
AOI22_X1 i_2348 (.ZN (n_2598), .A1 (inputB[18]), .A2 (inputA[14]), .B1 (inputB[19]), .B2 (inputA[13]));
INV_X1 i_2347 (.ZN (n_2597), .A (n_2598));
NAND2_X1 i_2346 (.ZN (n_2596), .A1 (n_2599), .A2 (n_2597));
NAND2_X1 i_2345 (.ZN (n_2595), .A1 (inputB[20]), .A2 (inputA[12]));
INV_X1 i_2344 (.ZN (n_2594), .A (n_2595));
XNOR2_X1 i_2343 (.ZN (n_3674), .A (n_2596), .B (n_2594));
AOI22_X1 i_2342 (.ZN (n_2592), .A1 (inputB[24]), .A2 (inputA[8]), .B1 (inputB[25]), .B2 (inputA[7]));
INV_X1 i_2341 (.ZN (n_2591), .A (n_2592));
AND2_X1 i_2340 (.ZN (n_2590), .A1 (inputB[25]), .A2 (inputA[8]));
NAND3_X1 i_2339 (.ZN (n_2589), .A1 (inputB[24]), .A2 (inputA[7]), .A3 (n_2590));
NAND2_X1 i_2338 (.ZN (n_2588), .A1 (n_2591), .A2 (n_2589));
NAND2_X1 i_2337 (.ZN (n_2586), .A1 (inputB[26]), .A2 (inputA[6]));
XOR2_X1 i_2336 (.Z (n_3660), .A (n_2588), .B (n_2586));
NAND2_X1 i_2335 (.ZN (n_2585), .A1 (inputB[28]), .A2 (inputA[5]));
INV_X1 i_2334 (.ZN (n_2584), .A (n_2585));
NAND2_X1 i_2333 (.ZN (n_2583), .A1 (n_2760), .A2 (n_2584));
AOI22_X1 i_2332 (.ZN (n_2582), .A1 (inputB[27]), .A2 (inputA[5]), .B1 (inputB[28]), .B2 (inputA[4]));
INV_X1 i_2331 (.ZN (n_2581), .A (n_2582));
NAND2_X1 i_2330 (.ZN (n_2578), .A1 (n_2583), .A2 (n_2581));
NAND2_X1 i_2329 (.ZN (n_2577), .A1 (inputB[29]), .A2 (inputA[3]));
XOR2_X1 i_2328 (.Z (n_3653), .A (n_2578), .B (n_2577));
AOI21_X1 i_2327 (.ZN (n_2573), .A (n_3571), .B1 (n_3570), .B2 (n_2738));
INV_X1 i_2326 (.ZN (n_3574), .A (n_2573));
AOI21_X1 i_2325 (.ZN (n_2568), .A (n_2752), .B1 (n_2748), .B2 (n_2745));
XOR2_X1 i_2324 (.Z (n_3734), .A (n_3732), .B (n_2568));
AOI22_X1 i_2323 (.ZN (n_2567), .A1 (n_2872), .A2 (n_2780), .B1 (n_2778), .B2 (n_2774));
XOR2_X1 i_2322 (.Z (n_3724), .A (n_3722), .B (n_2567));
AOI21_X1 i_2321 (.ZN (n_2563), .A (n_3586), .B1 (n_3585), .B2 (n_2679));
INV_X1 i_2320 (.ZN (n_3589), .A (n_2563));
AOI21_X1 i_2319 (.ZN (n_2559), .A (n_3576), .B1 (n_3575), .B2 (n_2719));
INV_X1 i_2318 (.ZN (n_3579), .A (n_2559));
AOI21_X1 i_2317 (.ZN (n_2558), .A (n_3591), .B1 (n_3590), .B2 (n_2733));
INV_X1 i_2316 (.ZN (n_3594), .A (n_2558));
AOI21_X1 i_2315 (.ZN (n_2557), .A (n_3601), .B1 (n_3600), .B2 (n_2714));
INV_X1 i_2314 (.ZN (n_3604), .A (n_2557));
AOI21_X1 i_2313 (.ZN (n_2553), .A (n_3596), .B1 (n_3595), .B2 (n_2673));
INV_X1 i_2312 (.ZN (n_3599), .A (n_2553));
NAND2_X1 i_2311 (.ZN (n_2548), .A1 (inputB[22]), .A2 (inputA[11]));
INV_X1 i_2310 (.ZN (n_2547), .A (n_2548));
NAND2_X1 i_2309 (.ZN (n_2543), .A1 (n_2766), .A2 (n_2547));
AOI22_X1 i_2308 (.ZN (n_2539), .A1 (inputB[21]), .A2 (inputA[11]), .B1 (inputB[22]), .B2 (inputA[10]));
INV_X1 i_2307 (.ZN (n_2538), .A (n_2539));
NAND2_X1 i_2306 (.ZN (n_2533), .A1 (n_2543), .A2 (n_2538));
NAND2_X1 i_2305 (.ZN (n_2528), .A1 (inputB[23]), .A2 (inputA[9]));
XOR2_X1 i_2304 (.Z (n_2527), .A (n_2533), .B (n_2528));
XOR2_X1 i_2303 (.Z (n_3754), .A (n_3752), .B (n_2527));
NAND2_X1 i_2302 (.ZN (n_2524), .A1 (inputB[13]), .A2 (inputA[20]));
INV_X1 i_2301 (.ZN (n_2523), .A (n_2524));
NAND2_X1 i_2300 (.ZN (n_2522), .A1 (n_2779), .A2 (n_2523));
AOI22_X1 i_2299 (.ZN (n_2518), .A1 (inputB[12]), .A2 (inputA[20]), .B1 (inputB[13]), .B2 (inputA[19]));
INV_X1 i_2297 (.ZN (n_2517), .A (n_2518));
NAND2_X1 i_2296 (.ZN (n_2514), .A1 (n_2522), .A2 (n_2517));
NAND2_X1 i_2295 (.ZN (n_2513), .A1 (inputB[14]), .A2 (inputA[18]));
XOR2_X1 i_2293 (.Z (n_2509), .A (n_2514), .B (n_2513));
XOR2_X1 i_2292 (.Z (n_3749), .A (n_3747), .B (n_2509));
AOI21_X1 i_2291 (.ZN (n_2508), .A (n_3606), .B1 (n_3605), .B2 (n_2704));
INV_X1 i_2289 (.ZN (n_3609), .A (n_2508));
AOI21_X1 i_2288 (.ZN (n_2507), .A (n_3581), .B1 (n_3580), .B2 (n_2726));
INV_X1 i_2287 (.ZN (n_2506), .A (n_2507));
XNOR2_X1 i_2285 (.ZN (n_3769), .A (n_3767), .B (n_2507));
AOI21_X1 i_2284 (.ZN (n_2503), .A (n_3611), .B1 (n_3610), .B2 (n_2675));
INV_X1 i_2283 (.ZN (n_3614), .A (n_2503));
AOI21_X1 i_2281 (.ZN (n_2502), .A (n_3556), .B1 (n_3555), .B2 (n_2674));
INV_X1 i_2280 (.ZN (n_2501), .A (n_2502));
XNOR2_X1 i_2279 (.ZN (n_2500), .A (n_3737), .B (n_2502));
XOR2_X1 i_2277 (.Z (n_3774), .A (n_3772), .B (n_2500));
AND2_X1 i_2276 (.ZN (n_2499), .A1 (inputB[31]), .A2 (inputA[1]));
NAND2_X1 i_2275 (.ZN (n_3649), .A1 (n_2749), .A2 (n_2499));
OAI21_X1 i_2273 (.ZN (n_2498), .A (n_3649), .B1 (n_2749), .B2 (n_2499));
XOR2_X1 i_2272 (.Z (n_2497), .A (n_3757), .B (n_2498));
XOR2_X1 i_2271 (.Z (n_3779), .A (n_3777), .B (n_2497));
AOI21_X1 i_2269 (.ZN (n_2496), .A (n_3621), .B1 (n_3620), .B2 (n_2669));
INV_X1 i_2268 (.ZN (n_3624), .A (n_2496));
AOI21_X1 i_2267 (.ZN (n_2495), .A (n_3626), .B1 (n_3625), .B2 (n_2650));
INV_X1 i_2265 (.ZN (n_3629), .A (n_2495));
NAND2_X1 i_2264 (.ZN (n_2494), .A1 (n_2763), .A2 (n_2761));
NAND2_X1 i_2263 (.ZN (n_2493), .A1 (n_2765), .A2 (n_2494));
XOR2_X1 i_2261 (.Z (n_2492), .A (n_3727), .B (n_2493));
XOR2_X1 i_2260 (.Z (n_2489), .A (n_3762), .B (n_2492));
XOR2_X1 i_2259 (.Z (n_3789), .A (n_3787), .B (n_2489));
AOI21_X1 i_2257 (.ZN (n_2488), .A (n_3631), .B1 (n_3630), .B2 (n_2658));
INV_X1 i_2256 (.ZN (n_3634), .A (n_2488));
NAND2_X1 i_2255 (.ZN (n_2487), .A1 (inputB[4]), .A2 (inputA[29]));
NAND2_X1 i_2253 (.ZN (n_2486), .A1 (inputB[4]), .A2 (inputA[28]));
OAI21_X1 i_2252 (.ZN (n_2485), .A (n_2486), .B1 (n_5756), .B2 (n_5750));
OAI21_X1 i_2251 (.ZN (n_2482), .A (n_2485), .B1 (n_2819), .B2 (n_2487));
NAND2_X1 i_2249 (.ZN (n_2481), .A1 (inputB[5]), .A2 (inputA[27]));
INV_X1 i_2248 (.ZN (n_2480), .A (n_2481));
XOR2_X1 i_2247 (.Z (n_2479), .A (n_2482), .B (n_2481));
XOR2_X1 i_2245 (.Z (n_2478), .A (n_3742), .B (n_2479));
XOR2_X1 i_2244 (.Z (n_2477), .A (n_3782), .B (n_2478));
XOR2_X1 i_2243 (.Z (n_3799), .A (n_3797), .B (n_2477));
AOI21_X1 i_2242 (.ZN (n_2476), .A (n_3616), .B1 (n_3615), .B2 (n_2699));
INV_X1 i_2241 (.ZN (n_2475), .A (n_2476));
XNOR2_X1 i_2240 (.ZN (n_2474), .A (n_3792), .B (n_2476));
XOR2_X1 i_2239 (.Z (n_3804), .A (n_3802), .B (n_2474));
AOI21_X1 i_2238 (.ZN (n_2473), .A (n_3636), .B1 (n_3635), .B2 (n_2649));
INV_X1 i_2237 (.ZN (n_2472), .A (n_2473));
XNOR2_X1 i_2236 (.ZN (n_3809), .A (n_3807), .B (n_2473));
NAND2_X1 i_2235 (.ZN (n_2471), .A1 (n_2485), .A2 (n_2480));
OAI21_X1 i_2234 (.ZN (n_3710), .A (n_2471), .B1 (n_2819), .B2 (n_2487));
OAI21_X1 i_2233 (.ZN (n_3703), .A (n_2623), .B1 (n_2627), .B2 (n_2619));
OAI21_X1 i_2232 (.ZN (n_3689), .A (n_2522), .B1 (n_2518), .B2 (n_2513));
OAI21_X1 i_2231 (.ZN (n_3682), .A (n_2606), .B1 (n_2611), .B2 (n_2609));
OAI21_X1 i_2230 (.ZN (n_3668), .A (n_2543), .B1 (n_2539), .B2 (n_2528));
OAI21_X1 i_2229 (.ZN (n_3661), .A (n_2589), .B1 (n_2592), .B2 (n_2586));
AOI21_X1 i_2228 (.ZN (n_2468), .A (n_3733), .B1 (n_3732), .B2 (n_2568));
INV_X1 i_2227 (.ZN (n_3736), .A (n_2468));
AOI21_X1 i_2226 (.ZN (n_2467), .A (n_3723), .B1 (n_3722), .B2 (n_2567));
INV_X1 i_2225 (.ZN (n_3726), .A (n_2467));
AND2_X1 i_2224 (.ZN (n_3717), .A1 (n_2638), .A2 (n_2631));
NAND2_X1 i_2223 (.ZN (n_2466), .A1 (inputB[6]), .A2 (inputA[28]));
INV_X1 i_2222 (.ZN (n_2465), .A (n_2466));
AOI22_X1 i_2221 (.ZN (n_2464), .A1 (inputB[5]), .A2 (inputA[28]), .B1 (inputB[6]), .B2 (inputA[27]));
AOI21_X1 i_2220 (.ZN (n_2461), .A (n_2464), .B1 (n_2480), .B2 (n_2465));
XOR2_X1 i_2219 (.Z (n_3876), .A (n_2624), .B (n_2461));
NAND2_X1 i_2218 (.ZN (n_2460), .A1 (inputB[9]), .A2 (inputA[25]));
NOR2_X1 i_2217 (.ZN (n_2459), .A1 (n_2619), .A2 (n_2460));
AOI22_X1 i_2216 (.ZN (n_2458), .A1 (inputB[8]), .A2 (inputA[25]), .B1 (inputB[9]), .B2 (inputA[24]));
NOR2_X1 i_2215 (.ZN (n_2457), .A1 (n_2459), .A2 (n_2458));
XOR2_X1 i_2214 (.Z (n_3869), .A (n_2618), .B (n_2457));
NAND2_X1 i_2213 (.ZN (n_2456), .A1 (inputB[15]), .A2 (inputA[19]));
NOR2_X1 i_2212 (.ZN (n_2455), .A1 (n_2513), .A2 (n_2456));
AOI22_X1 i_2211 (.ZN (n_2454), .A1 (inputB[14]), .A2 (inputA[19]), .B1 (inputB[15]), .B2 (inputA[18]));
NOR2_X1 i_2210 (.ZN (n_2453), .A1 (n_2455), .A2 (n_2454));
XOR2_X1 i_2209 (.Z (n_3855), .A (n_2607), .B (n_2453));
AOI22_X1 i_2208 (.ZN (n_2452), .A1 (inputB[17]), .A2 (inputA[16]), .B1 (inputB[18]), .B2 (inputA[15]));
INV_X1 i_2207 (.ZN (n_2451), .A (n_2452));
NAND3_X1 i_2206 (.ZN (n_2450), .A1 (inputB[18]), .A2 (inputA[16]), .A3 (n_2610));
NAND2_X1 i_2205 (.ZN (n_2447), .A1 (n_2451), .A2 (n_2450));
XNOR2_X1 i_2204 (.ZN (n_3848), .A (n_2602), .B (n_2447));
NAND2_X1 i_2203 (.ZN (n_2446), .A1 (inputB[24]), .A2 (inputA[10]));
NOR2_X1 i_2202 (.ZN (n_2442), .A1 (n_2528), .A2 (n_2446));
AOI22_X1 i_2201 (.ZN (n_2437), .A1 (inputB[23]), .A2 (inputA[10]), .B1 (inputB[24]), .B2 (inputA[9]));
NOR2_X1 i_2200 (.ZN (n_2436), .A1 (n_2442), .A2 (n_2437));
XOR2_X1 i_2199 (.Z (n_3834), .A (n_2590), .B (n_2436));
AOI22_X1 i_2198 (.ZN (n_2432), .A1 (inputB[26]), .A2 (inputA[7]), .B1 (inputB[27]), .B2 (inputA[6]));
INV_X1 i_2197 (.ZN (n_2428), .A (n_2432));
NAND4_X1 i_2196 (.ZN (n_2427), .A1 (inputB[26]), .A2 (inputA[7]), .A3 (inputB[27]), .A4 (inputA[6]));
NAND2_X1 i_2195 (.ZN (n_2426), .A1 (n_2428), .A2 (n_2427));
XNOR2_X1 i_2194 (.ZN (n_3827), .A (n_2584), .B (n_2426));
AOI21_X1 i_2193 (.ZN (n_2422), .A (n_3738), .B1 (n_3737), .B2 (n_2501));
INV_X1 i_2192 (.ZN (n_3741), .A (n_2422));
OAI21_X1 i_2191 (.ZN (n_2417), .A (n_2583), .B1 (n_2582), .B2 (n_2577));
XOR2_X1 i_2190 (.Z (n_3901), .A (n_3899), .B (n_2417));
OAI21_X1 i_2188 (.ZN (n_2412), .A (n_2617), .B1 (n_2616), .B2 (n_2612));
XOR2_X1 i_2187 (.Z (n_3891), .A (n_3889), .B (n_2412));
AOI21_X1 i_2186 (.ZN (n_2408), .A (n_3758), .B1 (n_3757), .B2 (n_2498));
INV_X1 i_2184 (.ZN (n_3761), .A (n_2408));
AOI21_X1 i_2183 (.ZN (n_2407), .A (n_3748), .B1 (n_3747), .B2 (n_2509));
INV_X1 i_2182 (.ZN (n_3751), .A (n_2407));
AOI21_X1 i_2180 (.ZN (n_2406), .A (n_3743), .B1 (n_3742), .B2 (n_2479));
INV_X1 i_2179 (.ZN (n_3746), .A (n_2406));
AOI21_X1 i_2178 (.ZN (n_2402), .A (n_3728), .B1 (n_3727), .B2 (n_2493));
INV_X1 i_2176 (.ZN (n_2397), .A (n_2402));
XNOR2_X1 i_2175 (.ZN (n_3906), .A (n_3904), .B (n_2402));
AOI21_X1 i_2174 (.ZN (n_2392), .A (n_3768), .B1 (n_3767), .B2 (n_2506));
INV_X1 i_2172 (.ZN (n_3771), .A (n_2392));
AOI22_X1 i_2171 (.ZN (n_2391), .A1 (inputB[29]), .A2 (inputA[4]), .B1 (inputB[30]), .B2 (inputA[3]));
INV_X1 i_2170 (.ZN (n_2387), .A (n_2391));
NAND4_X1 i_2168 (.ZN (n_2382), .A1 (inputB[29]), .A2 (inputA[3]), .A3 (inputB[30]), .A4 (inputA[4]));
NAND2_X1 i_2167 (.ZN (n_2378), .A1 (n_2387), .A2 (n_2382));
NAND2_X1 i_2166 (.ZN (n_2377), .A1 (inputB[31]), .A2 (inputA[2]));
INV_X1 i_2164 (.ZN (n_2376), .A (n_2377));
XNOR2_X1 i_2163 (.ZN (n_2375), .A (n_2378), .B (n_2377));
XOR2_X1 i_2162 (.Z (n_3926), .A (n_3924), .B (n_2375));
AND2_X1 i_2160 (.ZN (n_2373), .A1 (inputB[21]), .A2 (inputA[13]));
NAND2_X1 i_2159 (.ZN (n_2372), .A1 (n_2594), .A2 (n_2373));
AOI22_X1 i_2158 (.ZN (n_2371), .A1 (inputB[20]), .A2 (inputA[13]), .B1 (inputB[21]), .B2 (inputA[12]));
AOI21_X1 i_2156 (.ZN (n_2370), .A (n_2371), .B1 (n_2594), .B2 (n_2373));
XOR2_X1 i_2155 (.Z (n_2369), .A (n_2547), .B (n_2370));
XOR2_X1 i_2154 (.Z (n_3921), .A (n_3919), .B (n_2369));
AOI21_X1 i_2152 (.ZN (n_2368), .A (n_3773), .B1 (n_3772), .B2 (n_2500));
INV_X1 i_2151 (.ZN (n_3776), .A (n_2368));
AOI211_X1 i_2150 (.ZN (n_2367), .A (n_5755), .B (n_5753), .C1 (inputB[3]), .C2 (inputA[30]));
INV_X1 i_2148 (.ZN (n_2366), .A (n_2367));
OAI211_X1 i_2147 (.ZN (n_2365), .A (inputB[3]), .B (inputA[30]), .C1 (n_5755), .C2 (n_5753));
NAND2_X1 i_2146 (.ZN (n_2364), .A1 (n_2366), .A2 (n_2365));
XOR2_X1 i_2144 (.Z (n_2363), .A (n_2487), .B (n_2364));
XOR2_X1 i_2143 (.Z (n_2362), .A (n_3909), .B (n_2363));
XOR2_X1 i_2142 (.Z (n_3941), .A (n_3939), .B (n_2362));
AOI21_X1 i_2140 (.ZN (n_2359), .A (n_2598), .B1 (n_2599), .B2 (n_2595));
XOR2_X1 i_2139 (.Z (n_2358), .A (n_3894), .B (n_2359));
XOR2_X1 i_2138 (.Z (n_3931), .A (n_3929), .B (n_2358));
AOI21_X1 i_2137 (.ZN (n_2357), .A (n_3783), .B1 (n_3782), .B2 (n_2478));
INV_X1 i_2136 (.ZN (n_3786), .A (n_2357));
AOI21_X1 i_2135 (.ZN (n_2356), .A (n_3763), .B1 (n_3762), .B2 (n_2492));
INV_X1 i_2134 (.ZN (n_2355), .A (n_2356));
XNOR2_X1 i_2133 (.ZN (n_3946), .A (n_3944), .B (n_2356));
AOI21_X1 i_2132 (.ZN (n_2352), .A (n_3788), .B1 (n_3787), .B2 (n_2489));
INV_X1 i_2131 (.ZN (n_3791), .A (n_2352));
AND2_X1 i_2130 (.ZN (n_2351), .A1 (inputB[12]), .A2 (inputA[22]));
NAND3_X1 i_2129 (.ZN (n_2350), .A1 (inputB[11]), .A2 (inputA[21]), .A3 (n_2351));
AOI22_X1 i_2128 (.ZN (n_2349), .A1 (inputB[11]), .A2 (inputA[22]), .B1 (inputB[12]), .B2 (inputA[21]));
INV_X1 i_2127 (.ZN (n_2348), .A (n_2349));
NAND2_X1 i_2126 (.ZN (n_2347), .A1 (n_2350), .A2 (n_2348));
XNOR2_X1 i_2125 (.ZN (n_2346), .A (n_2523), .B (n_2347));
XOR2_X1 i_2124 (.Z (n_2345), .A (n_3914), .B (n_2346));
XOR2_X1 i_2123 (.Z (n_3951), .A (n_3949), .B (n_2345));
AOI21_X1 i_2122 (.ZN (n_2344), .A (n_3778), .B1 (n_3777), .B2 (n_2497));
INV_X1 i_2121 (.ZN (n_2343), .A (n_2344));
XNOR2_X1 i_2120 (.ZN (n_3961), .A (n_3959), .B (n_2344));
AOI21_X1 i_2119 (.ZN (n_2342), .A (n_3798), .B1 (n_3797), .B2 (n_2477));
INV_X1 i_2118 (.ZN (n_3801), .A (n_2342));
AOI21_X1 i_2117 (.ZN (n_2341), .A (n_3793), .B1 (n_3792), .B2 (n_2475));
INV_X1 i_2116 (.ZN (n_2338), .A (n_2341));
XNOR2_X1 i_2115 (.ZN (n_3966), .A (n_3964), .B (n_2341));
AOI21_X1 i_2114 (.ZN (n_2337), .A (n_3753), .B1 (n_3752), .B2 (n_2527));
INV_X1 i_2113 (.ZN (n_2336), .A (n_2337));
XNOR2_X1 i_2112 (.ZN (n_2335), .A (n_3934), .B (n_2337));
XOR2_X1 i_2111 (.Z (n_2334), .A (n_3954), .B (n_2335));
XOR2_X1 i_2110 (.Z (n_3971), .A (n_3969), .B (n_2334));
AOI21_X1 i_2109 (.ZN (n_2331), .A (n_3808), .B1 (n_3807), .B2 (n_2472));
INV_X1 i_2108 (.ZN (n_3811), .A (n_2331));
OAI22_X1 i_2107 (.ZN (n_3877), .A1 (n_2481), .A2 (n_2466), .B1 (n_2625), .B2 (n_2464));
NOR2_X1 i_2106 (.ZN (n_2330), .A1 (n_2618), .A2 (n_2459));
NOR2_X1 i_2105 (.ZN (n_3870), .A1 (n_2458), .A2 (n_2330));
NOR2_X1 i_2104 (.ZN (n_2329), .A1 (n_2607), .A2 (n_2455));
NOR2_X1 i_2103 (.ZN (n_3856), .A1 (n_2454), .A2 (n_2329));
OAI21_X1 i_2102 (.ZN (n_3849), .A (n_2450), .B1 (n_2603), .B2 (n_2452));
NOR2_X1 i_2101 (.ZN (n_2328), .A1 (n_2590), .A2 (n_2442));
NOR2_X1 i_2100 (.ZN (n_3835), .A1 (n_2437), .A2 (n_2328));
OAI21_X1 i_2099 (.ZN (n_3828), .A (n_2427), .B1 (n_2585), .B2 (n_2432));
AOI21_X1 i_2098 (.ZN (n_2327), .A (n_3900), .B1 (n_3899), .B2 (n_2417));
INV_X1 i_2097 (.ZN (n_3903), .A (n_2327));
AOI21_X1 i_2096 (.ZN (n_2326), .A (n_3895), .B1 (n_3894), .B2 (n_2359));
INV_X1 i_2095 (.ZN (n_3898), .A (n_2326));
AOI211_X1 i_2094 (.ZN (n_2325), .A (n_5756), .B (n_5753), .C1 (inputB[4]), .C2 (inputA[30]));
OAI211_X1 i_2093 (.ZN (n_2324), .A (inputB[4]), .B (inputA[30]), .C1 (n_5756), .C2 (n_5753));
INV_X1 i_2092 (.ZN (n_2323), .A (n_2324));
NOR2_X1 i_2091 (.ZN (n_2319), .A1 (n_2325), .A2 (n_2323));
AOI21_X1 i_2090 (.ZN (n_2314), .A (n_2367), .B1 (n_2487), .B2 (n_2365));
INV_X1 i_2089 (.ZN (n_2313), .A (n_2314));
XOR2_X1 i_2088 (.Z (n_4050), .A (n_2319), .B (n_2314));
NAND2_X1 i_2087 (.ZN (n_2309), .A1 (inputB[5]), .A2 (inputA[29]));
NOR2_X1 i_2086 (.ZN (n_2305), .A1 (n_2466), .A2 (n_2309));
INV_X1 i_2085 (.ZN (n_2304), .A (n_2305));
AOI21_X1 i_2084 (.ZN (n_2303), .A (n_2305), .B1 (n_2466), .B2 (n_2309));
NAND2_X1 i_2082 (.ZN (n_2300), .A1 (inputB[7]), .A2 (inputA[27]));
XNOR2_X1 i_2081 (.ZN (n_4043), .A (n_2303), .B (n_2300));
AOI21_X1 i_2080 (.ZN (n_2299), .A (n_2351), .B1 (inputB[11]), .B2 (inputA[23]));
INV_X1 i_2078 (.ZN (n_2294), .A (n_2299));
NAND3_X1 i_2077 (.ZN (n_2289), .A1 (inputB[11]), .A2 (inputA[23]), .A3 (n_2351));
NAND2_X1 i_2076 (.ZN (n_2288), .A1 (n_2294), .A2 (n_2289));
NAND2_X1 i_2074 (.ZN (n_2285), .A1 (inputB[13]), .A2 (inputA[21]));
XOR2_X1 i_2073 (.Z (n_4029), .A (n_2288), .B (n_2285));
NAND2_X1 i_2072 (.ZN (n_2284), .A1 (inputB[14]), .A2 (inputA[20]));
NOR2_X1 i_2070 (.ZN (n_2279), .A1 (n_2456), .A2 (n_2284));
AOI21_X1 i_2069 (.ZN (n_2274), .A (n_2279), .B1 (n_2456), .B2 (n_2284));
AND2_X1 i_2068 (.ZN (n_2269), .A1 (inputB[16]), .A2 (inputA[18]));
XOR2_X1 i_2066 (.Z (n_4022), .A (n_2274), .B (n_2269));
AOI21_X1 i_2065 (.ZN (n_2268), .A (n_2373), .B1 (inputB[20]), .B2 (inputA[14]));
INV_X1 i_2064 (.ZN (n_2265), .A (n_2268));
NAND3_X1 i_2062 (.ZN (n_2264), .A1 (inputB[20]), .A2 (inputA[14]), .A3 (n_2373));
NAND2_X1 i_2061 (.ZN (n_2260), .A1 (n_2265), .A2 (n_2264));
NAND2_X1 i_2060 (.ZN (n_2259), .A1 (inputB[22]), .A2 (inputA[12]));
XOR2_X1 i_2058 (.Z (n_4008), .A (n_2260), .B (n_2259));
NAND2_X1 i_2057 (.ZN (n_2258), .A1 (inputB[23]), .A2 (inputA[11]));
NOR2_X1 i_2056 (.ZN (n_2257), .A1 (n_2446), .A2 (n_2258));
INV_X1 i_2054 (.ZN (n_2256), .A (n_2257));
AOI21_X1 i_2053 (.ZN (n_2254), .A (n_2257), .B1 (n_2446), .B2 (n_2258));
NAND2_X1 i_2052 (.ZN (n_2253), .A1 (inputB[25]), .A2 (inputA[9]));
XNOR2_X1 i_2050 (.ZN (n_4001), .A (n_2254), .B (n_2253));
AND2_X1 i_2049 (.ZN (n_2252), .A1 (inputB[31]), .A2 (inputA[3]));
AOI22_X1 i_2048 (.ZN (n_2251), .A1 (inputB[30]), .A2 (inputA[4]), .B1 (inputB[29]), .B2 (inputA[5]));
INV_X1 i_2046 (.ZN (n_2250), .A (n_2251));
NAND2_X1 i_2045 (.ZN (n_2247), .A1 (inputB[30]), .A2 (inputA[5]));
INV_X1 i_2044 (.ZN (n_2246), .A (n_2247));
NAND3_X1 i_2042 (.ZN (n_2245), .A1 (inputB[29]), .A2 (inputA[4]), .A3 (n_2246));
NAND2_X1 i_2041 (.ZN (n_2244), .A1 (n_2250), .A2 (n_2245));
XOR2_X1 i_2040 (.Z (n_3985), .A (n_2252), .B (n_2244));
AOI21_X1 i_2038 (.ZN (n_2243), .A (n_3905), .B1 (n_3904), .B2 (n_2397));
INV_X1 i_2037 (.ZN (n_3908), .A (n_2243));
OAI21_X1 i_2036 (.ZN (n_2240), .A (n_2372), .B1 (n_2548), .B2 (n_2371));
XOR2_X1 i_2035 (.Z (n_4063), .A (n_4061), .B (n_2240));
AOI21_X1 i_2034 (.ZN (n_2239), .A (n_2349), .B1 (n_2524), .B2 (n_2350));
XOR2_X1 i_2033 (.Z (n_4058), .A (n_4056), .B (n_2239));
AOI21_X1 i_2032 (.ZN (n_2238), .A (n_3920), .B1 (n_3919), .B2 (n_2369));
INV_X1 i_2031 (.ZN (n_3923), .A (n_2238));
AOI21_X1 i_2030 (.ZN (n_2237), .A (n_3915), .B1 (n_3914), .B2 (n_2346));
INV_X1 i_2029 (.ZN (n_3918), .A (n_2237));
AOI21_X1 i_2028 (.ZN (n_2236), .A (n_3890), .B1 (n_3889), .B2 (n_2412));
INV_X1 i_2027 (.ZN (n_2235), .A (n_2236));
XNOR2_X1 i_2026 (.ZN (n_4073), .A (n_4071), .B (n_2236));
AOI21_X1 i_2025 (.ZN (n_2234), .A (n_3935), .B1 (n_3934), .B2 (n_2336));
INV_X1 i_2024 (.ZN (n_3938), .A (n_2234));
NAND2_X1 i_2023 (.ZN (n_2233), .A1 (inputB[27]), .A2 (inputA[8]));
INV_X1 i_2022 (.ZN (n_2232), .A (n_2233));
NAND3_X1 i_2021 (.ZN (n_2231), .A1 (inputB[26]), .A2 (inputA[7]), .A3 (n_2232));
AOI22_X1 i_2020 (.ZN (n_2230), .A1 (inputB[27]), .A2 (inputA[7]), .B1 (inputB[26]), .B2 (inputA[8]));
INV_X1 i_2019 (.ZN (n_2229), .A (n_2230));
NAND2_X1 i_2018 (.ZN (n_2226), .A1 (n_2231), .A2 (n_2229));
NAND2_X1 i_2017 (.ZN (n_2225), .A1 (inputB[28]), .A2 (inputA[6]));
XOR2_X1 i_2016 (.Z (n_2224), .A (n_2226), .B (n_2225));
XOR2_X1 i_2015 (.Z (n_4088), .A (n_4086), .B (n_2224));
AND2_X1 i_2014 (.ZN (n_2223), .A1 (inputB[18]), .A2 (inputA[17]));
NAND3_X1 i_2013 (.ZN (n_2222), .A1 (inputB[17]), .A2 (inputA[16]), .A3 (n_2223));
AOI22_X1 i_2012 (.ZN (n_2219), .A1 (inputB[18]), .A2 (inputA[16]), .B1 (inputB[17]), .B2 (inputA[17]));
INV_X1 i_2011 (.ZN (n_2218), .A (n_2219));
NAND2_X1 i_2010 (.ZN (n_2217), .A1 (n_2222), .A2 (n_2218));
NAND2_X1 i_2009 (.ZN (n_2216), .A1 (inputB[19]), .A2 (inputA[15]));
XOR2_X1 i_2008 (.Z (n_2215), .A (n_2217), .B (n_2216));
XOR2_X1 i_2007 (.Z (n_4083), .A (n_4081), .B (n_2215));
AOI21_X1 i_2006 (.ZN (n_2214), .A (n_2391), .B1 (n_2382), .B2 (n_2376));
XOR2_X1 i_2005 (.Z (n_2213), .A (n_4066), .B (n_2214));
XOR2_X1 i_2004 (.Z (n_4093), .A (n_4091), .B (n_2213));
AOI21_X1 i_2003 (.ZN (n_2212), .A (n_3945), .B1 (n_3944), .B2 (n_2355));
INV_X1 i_2002 (.ZN (n_3948), .A (n_2212));
AOI21_X1 i_2001 (.ZN (n_2211), .A (n_3910), .B1 (n_3909), .B2 (n_2363));
INV_X1 i_2000 (.ZN (n_2210), .A (n_2211));
XNOR2_X1 i_1999 (.ZN (n_4103), .A (n_4101), .B (n_2211));
AOI21_X1 i_1998 (.ZN (n_2209), .A (n_3925), .B1 (n_3924), .B2 (n_2375));
INV_X1 i_1997 (.ZN (n_2208), .A (n_2209));
XNOR2_X1 i_1996 (.ZN (n_4098), .A (n_4096), .B (n_2209));
AOI21_X1 i_1995 (.ZN (n_2205), .A (n_3930), .B1 (n_3929), .B2 (n_2358));
INV_X1 i_1994 (.ZN (n_2204), .A (n_2205));
XNOR2_X1 i_1993 (.ZN (n_4108), .A (n_4106), .B (n_2205));
AOI21_X1 i_1992 (.ZN (n_2200), .A (n_3960), .B1 (n_3959), .B2 (n_2343));
INV_X1 i_1991 (.ZN (n_3963), .A (n_2200));
NAND2_X1 i_1990 (.ZN (n_2195), .A1 (inputB[8]), .A2 (inputA[26]));
NAND2_X1 i_1989 (.ZN (n_2194), .A1 (n_2460), .A2 (n_2195));
INV_X1 i_1988 (.ZN (n_2190), .A (n_2194));
OAI21_X1 i_1987 (.ZN (n_2186), .A (n_2194), .B1 (n_2460), .B2 (n_2195));
NAND2_X1 i_1986 (.ZN (n_2185), .A1 (inputB[10]), .A2 (inputA[24]));
XOR2_X1 i_1985 (.Z (n_2184), .A (n_2186), .B (n_2185));
XOR2_X1 i_1984 (.Z (n_2180), .A (n_4076), .B (n_2184));
XOR2_X1 i_1983 (.Z (n_4113), .A (n_4111), .B (n_2180));
AOI21_X1 i_1982 (.ZN (n_2175), .A (n_3940), .B1 (n_3939), .B2 (n_2362));
INV_X1 i_1980 (.ZN (n_2174), .A (n_2175));
XNOR2_X1 i_1979 (.ZN (n_4118), .A (n_4116), .B (n_2175));
AOI21_X1 i_1978 (.ZN (n_2171), .A (n_3950), .B1 (n_3949), .B2 (n_2345));
INV_X1 i_1976 (.ZN (n_2170), .A (n_2171));
XNOR2_X1 i_1975 (.ZN (n_4123), .A (n_4121), .B (n_2171));
AOI21_X1 i_1974 (.ZN (n_2165), .A (n_3955), .B1 (n_3954), .B2 (n_2335));
INV_X1 i_1972 (.ZN (n_2161), .A (n_2165));
XNOR2_X1 i_1971 (.ZN (n_4128), .A (n_4126), .B (n_2165));
AOI21_X1 i_1970 (.ZN (n_2160), .A (n_3965), .B1 (n_3964), .B2 (n_2338));
INV_X1 i_1968 (.ZN (n_2159), .A (n_2160));
XNOR2_X1 i_1967 (.ZN (n_4133), .A (n_4131), .B (n_2160));
AOI21_X1 i_1966 (.ZN (n_2155), .A (n_3803), .B1 (n_3802), .B2 (n_2474));
INV_X1 i_1964 (.ZN (n_2154), .A (n_2155));
AOI21_X1 i_1963 (.ZN (n_2150), .A (n_3975), .B1 (n_3974), .B2 (n_2154));
INV_X1 i_1962 (.ZN (n_3978), .A (n_2150));
NAND2_X1 i_1960 (.ZN (n_384), .A1 (inputB[4]), .A2 (inputA[31]));
AOI22_X1 i_1959 (.ZN (n_4044), .A1 (n_2466), .A2 (n_2309), .B1 (n_2304), .B2 (n_2300));
OAI21_X1 i_1958 (.ZN (n_4030), .A (n_2289), .B1 (n_2299), .B2 (n_2285));
NOR2_X1 i_1956 (.ZN (n_2146), .A1 (n_2279), .A2 (n_2269));
AOI21_X1 i_1955 (.ZN (n_4023), .A (n_2146), .B1 (n_2456), .B2 (n_2284));
OAI21_X1 i_1954 (.ZN (n_4009), .A (n_2264), .B1 (n_2268), .B2 (n_2259));
AOI22_X1 i_1952 (.ZN (n_4002), .A1 (n_2446), .A2 (n_2258), .B1 (n_2256), .B2 (n_2253));
OAI21_X1 i_1951 (.ZN (n_3986), .A (n_2245), .B1 (n_2252), .B2 (n_2251));
AOI21_X1 i_1950 (.ZN (n_2145), .A (n_4067), .B1 (n_4066), .B2 (n_2214));
INV_X1 i_1948 (.ZN (n_4070), .A (n_2145));
AOI21_X1 i_1947 (.ZN (n_2144), .A (n_4057), .B1 (n_4056), .B2 (n_2239));
INV_X1 i_1946 (.ZN (n_4060), .A (n_2144));
AOI21_X1 i_1944 (.ZN (n_4051), .A (n_2325), .B1 (n_2324), .B2 (n_2313));
AOI22_X1 i_1943 (.ZN (n_2143), .A1 (inputB[9]), .A2 (inputA[26]), .B1 (inputB[8]), .B2 (inputA[27]));
INV_X1 i_1942 (.ZN (n_2140), .A (n_2143));
NAND4_X1 i_1940 (.ZN (n_2139), .A1 (inputB[8]), .A2 (inputA[26]), .A3 (inputB[9]), .A4 (inputA[27]));
NAND2_X1 i_1939 (.ZN (n_2138), .A1 (n_2140), .A2 (n_2139));
NAND2_X1 i_1938 (.ZN (n_2137), .A1 (inputB[10]), .A2 (inputA[25]));
XOR2_X1 i_1936 (.Z (n_4198), .A (n_2138), .B (n_2137));
AND2_X1 i_1935 (.ZN (n_2136), .A1 (inputB[11]), .A2 (inputA[24]));
AOI21_X1 i_1934 (.ZN (n_2135), .A (n_2136), .B1 (inputB[12]), .B2 (inputA[23]));
INV_X1 i_1933 (.ZN (n_2133), .A (n_2135));
NAND3_X1 i_1932 (.ZN (n_2132), .A1 (inputB[12]), .A2 (inputA[23]), .A3 (n_2136));
NAND2_X1 i_1931 (.ZN (n_2131), .A1 (n_2133), .A2 (n_2132));
NAND2_X1 i_1930 (.ZN (n_2130), .A1 (inputB[13]), .A2 (inputA[22]));
XOR2_X1 i_1929 (.Z (n_4191), .A (n_2131), .B (n_2130));
AOI21_X1 i_1928 (.ZN (n_2129), .A (n_2223), .B1 (inputB[17]), .B2 (inputA[18]));
INV_X1 i_1927 (.ZN (n_2127), .A (n_2129));
NAND3_X1 i_1926 (.ZN (n_2126), .A1 (inputB[17]), .A2 (inputA[18]), .A3 (n_2223));
NAND2_X1 i_1925 (.ZN (n_2125), .A1 (n_2127), .A2 (n_2126));
NAND2_X1 i_1924 (.ZN (n_2124), .A1 (inputB[19]), .A2 (inputA[16]));
XOR2_X1 i_1923 (.Z (n_4177), .A (n_2125), .B (n_2124));
AND2_X1 i_1922 (.ZN (n_2123), .A1 (inputB[20]), .A2 (inputA[15]));
AOI21_X1 i_1921 (.ZN (n_2122), .A (n_2123), .B1 (inputB[21]), .B2 (inputA[14]));
INV_X1 i_1920 (.ZN (n_2119), .A (n_2122));
NAND3_X1 i_1919 (.ZN (n_2118), .A1 (inputB[21]), .A2 (inputA[14]), .A3 (n_2123));
NAND2_X1 i_1918 (.ZN (n_2117), .A1 (n_2119), .A2 (n_2118));
NAND2_X1 i_1917 (.ZN (n_2116), .A1 (inputB[22]), .A2 (inputA[13]));
XOR2_X1 i_1916 (.Z (n_4170), .A (n_2117), .B (n_2116));
NAND2_X1 i_1915 (.ZN (n_2115), .A1 (inputB[26]), .A2 (inputA[9]));
INV_X1 i_1914 (.ZN (n_2114), .A (n_2115));
NAND2_X1 i_1913 (.ZN (n_2112), .A1 (n_2232), .A2 (n_2114));
OAI21_X1 i_1912 (.ZN (n_2111), .A (n_2112), .B1 (n_2232), .B2 (n_2114));
NAND2_X1 i_1911 (.ZN (n_2110), .A1 (inputB[28]), .A2 (inputA[7]));
XOR2_X1 i_1910 (.Z (n_4156), .A (n_2111), .B (n_2110));
NAND2_X1 i_1909 (.ZN (n_2109), .A1 (inputB[29]), .A2 (inputA[6]));
INV_X1 i_1908 (.ZN (n_2108), .A (n_2109));
NAND2_X1 i_1907 (.ZN (n_2106), .A1 (n_2246), .A2 (n_2108));
NAND2_X1 i_1906 (.ZN (n_2105), .A1 (n_2247), .A2 (n_2109));
AND2_X1 i_1905 (.ZN (n_2104), .A1 (n_2106), .A2 (n_2105));
NAND2_X1 i_1904 (.ZN (n_2103), .A1 (inputB[31]), .A2 (inputA[4]));
XOR2_X1 i_1903 (.Z (n_4147), .A (n_2104), .B (n_2103));
AOI21_X1 i_1902 (.ZN (n_2102), .A (n_2230), .B1 (n_2231), .B2 (n_2225));
XOR2_X1 i_1901 (.Z (n_4222), .A (n_4220), .B (n_2102));
AOI21_X1 i_1900 (.ZN (n_2101), .A (n_2219), .B1 (n_2222), .B2 (n_2216));
XOR2_X1 i_1899 (.Z (n_4217), .A (n_4215), .B (n_2101));
AOI21_X1 i_1898 (.ZN (n_2098), .A (n_4087), .B1 (n_4086), .B2 (n_2224));
INV_X1 i_1897 (.ZN (n_4090), .A (n_2098));
AOI21_X1 i_1896 (.ZN (n_2097), .A (n_4082), .B1 (n_4081), .B2 (n_2215));
INV_X1 i_1895 (.ZN (n_4085), .A (n_2097));
NAND2_X1 i_1894 (.ZN (n_2096), .A1 (inputB[6]), .A2 (inputA[30]));
OR2_X1 i_1893 (.ZN (n_2095), .A1 (n_2309), .A2 (n_2096));
AOI22_X1 i_1892 (.ZN (n_2094), .A1 (inputB[6]), .A2 (inputA[29]), .B1 (inputB[5]), .B2 (inputA[30]));
INV_X1 i_1891 (.ZN (n_2093), .A (n_2094));
NAND2_X1 i_1890 (.ZN (n_2091), .A1 (n_2095), .A2 (n_2093));
NAND2_X1 i_1889 (.ZN (n_2090), .A1 (inputB[7]), .A2 (inputA[28]));
XOR2_X1 i_1888 (.Z (n_2086), .A (n_2091), .B (n_2090));
XOR2_X1 i_1886 (.Z (n_4232), .A (n_4230), .B (n_2086));
AOI21_X1 i_1885 (.ZN (n_2081), .A (n_4062), .B1 (n_4061), .B2 (n_2240));
INV_X1 i_1884 (.ZN (n_2080), .A (n_2081));
XNOR2_X1 i_1882 (.ZN (n_4227), .A (n_4225), .B (n_2081));
AOI21_X1 i_1881 (.ZN (n_2076), .A (n_4097), .B1 (n_4096), .B2 (n_2208));
INV_X1 i_1880 (.ZN (n_4100), .A (n_2076));
AOI21_X1 i_1878 (.ZN (n_2071), .A (n_4092), .B1 (n_4091), .B2 (n_2213));
INV_X1 i_1877 (.ZN (n_4095), .A (n_2071));
NAND2_X1 i_1876 (.ZN (n_2070), .A1 (inputB[24]), .A2 (inputA[12]));
AOI22_X1 i_1874 (.ZN (n_2066), .A1 (inputB[24]), .A2 (inputA[11]), .B1 (inputB[23]), .B2 (inputA[12]));
INV_X1 i_1873 (.ZN (n_2062), .A (n_2066));
OAI21_X1 i_1872 (.ZN (n_2061), .A (n_2062), .B1 (n_2258), .B2 (n_2070));
NAND2_X1 i_1870 (.ZN (n_2060), .A1 (inputB[25]), .A2 (inputA[10]));
XOR2_X1 i_1869 (.Z (n_2057), .A (n_2061), .B (n_2060));
XOR2_X1 i_1868 (.Z (n_4242), .A (n_4240), .B (n_2057));
NAND2_X1 i_1866 (.ZN (n_2056), .A1 (inputB[15]), .A2 (inputA[21]));
AOI22_X1 i_1865 (.ZN (n_2055), .A1 (inputB[15]), .A2 (inputA[20]), .B1 (inputB[14]), .B2 (inputA[21]));
INV_X1 i_1864 (.ZN (n_2051), .A (n_2055));
OAI21_X1 i_1862 (.ZN (n_2046), .A (n_2051), .B1 (n_2284), .B2 (n_2056));
NAND2_X1 i_1861 (.ZN (n_2045), .A1 (inputB[16]), .A2 (inputA[19]));
XOR2_X1 i_1860 (.Z (n_2042), .A (n_2046), .B (n_2045));
XOR2_X1 i_1858 (.Z (n_4237), .A (n_4235), .B (n_2042));
AOI21_X1 i_1857 (.ZN (n_2041), .A (n_4077), .B1 (n_4076), .B2 (n_2184));
INV_X1 i_1856 (.ZN (n_2036), .A (n_2041));
XNOR2_X1 i_1854 (.ZN (n_4257), .A (n_4255), .B (n_2041));
OAI22_X1 i_1853 (.ZN (n_2035), .A1 (n_2460), .A2 (n_2195), .B1 (n_2190), .B2 (n_2185));
XOR2_X1 i_1852 (.Z (n_2032), .A (n_4210), .B (n_2035));
XOR2_X1 i_1850 (.Z (n_4252), .A (n_4250), .B (n_2032));
AOI21_X1 i_1849 (.ZN (n_2031), .A (n_4117), .B1 (n_4116), .B2 (n_2174));
INV_X1 i_1848 (.ZN (n_4120), .A (n_2031));
AOI21_X1 i_1846 (.ZN (n_2030), .A (n_4072), .B1 (n_4071), .B2 (n_2235));
INV_X1 i_1845 (.ZN (n_2029), .A (n_2030));
XNOR2_X1 i_1844 (.ZN (n_2028), .A (n_4245), .B (n_2030));
XOR2_X1 i_1843 (.Z (n_4267), .A (n_4265), .B (n_2028));
AOI21_X1 i_1842 (.ZN (n_2027), .A (n_4122), .B1 (n_4121), .B2 (n_2170));
INV_X1 i_1841 (.ZN (n_4125), .A (n_2027));
AOI21_X1 i_1840 (.ZN (n_2026), .A (n_4107), .B1 (n_4106), .B2 (n_2204));
INV_X1 i_1839 (.ZN (n_2025), .A (n_2026));
XNOR2_X1 i_1838 (.ZN (n_4272), .A (n_4270), .B (n_2026));
AOI21_X1 i_1837 (.ZN (n_2024), .A (n_4112), .B1 (n_4111), .B2 (n_2180));
INV_X1 i_1836 (.ZN (n_2023), .A (n_2024));
XNOR2_X1 i_1835 (.ZN (n_4277), .A (n_4275), .B (n_2024));
AOI21_X1 i_1834 (.ZN (n_2022), .A (n_4132), .B1 (n_4131), .B2 (n_2159));
INV_X1 i_1833 (.ZN (n_4135), .A (n_2022));
AOI21_X1 i_1832 (.ZN (n_2020), .A (n_4127), .B1 (n_4126), .B2 (n_2161));
INV_X1 i_1831 (.ZN (n_2019), .A (n_2020));
XNOR2_X1 i_1830 (.ZN (n_4287), .A (n_4285), .B (n_2020));
AOI21_X1 i_1829 (.ZN (n_2018), .A (n_3970), .B1 (n_3969), .B2 (n_2334));
INV_X1 i_1828 (.ZN (n_2017), .A (n_2018));
AOI21_X1 i_1827 (.ZN (n_2016), .A (n_4137), .B1 (n_4136), .B2 (n_2017));
INV_X1 i_1826 (.ZN (n_4140), .A (n_2016));
AOI21_X1 i_1825 (.ZN (n_4206), .A (n_2094), .B1 (n_2095), .B2 (n_2090));
OAI21_X1 i_1824 (.ZN (n_4199), .A (n_2139), .B1 (n_2143), .B2 (n_2137));
OAI22_X1 i_1823 (.ZN (n_4185), .A1 (n_2284), .A2 (n_2056), .B1 (n_2055), .B2 (n_2045));
OAI21_X1 i_1822 (.ZN (n_4178), .A (n_2126), .B1 (n_2129), .B2 (n_2124));
OAI22_X1 i_1821 (.ZN (n_4164), .A1 (n_2258), .A2 (n_2070), .B1 (n_2066), .B2 (n_2060));
AOI22_X1 i_1820 (.ZN (n_4157), .A1 (n_2233), .A2 (n_2115), .B1 (n_2112), .B2 (n_2110));
AOI21_X1 i_1819 (.ZN (n_2013), .A (n_4221), .B1 (n_4220), .B2 (n_2102));
INV_X1 i_1818 (.ZN (n_4224), .A (n_2013));
AOI21_X1 i_1817 (.ZN (n_2012), .A (n_4216), .B1 (n_4215), .B2 (n_2101));
INV_X1 i_1816 (.ZN (n_4219), .A (n_2012));
AOI21_X1 i_1815 (.ZN (n_2011), .A (n_2096), .B1 (inputB[5]), .B2 (inputA[31]));
INV_X1 i_1814 (.ZN (n_2010), .A (n_2011));
AND3_X1 i_1813 (.ZN (n_2009), .A1 (inputB[5]), .A2 (inputA[31]), .A3 (n_2096));
NOR2_X1 i_1812 (.ZN (n_2007), .A1 (n_2011), .A2 (n_2009));
NAND2_X1 i_1811 (.ZN (n_2006), .A1 (inputB[7]), .A2 (inputA[29]));
XNOR2_X1 i_1810 (.ZN (n_4358), .A (n_2007), .B (n_2006));
AOI22_X1 i_1809 (.ZN (n_2005), .A1 (inputB[9]), .A2 (inputA[27]), .B1 (inputB[8]), .B2 (inputA[28]));
INV_X1 i_1808 (.ZN (n_2004), .A (n_2005));
NAND2_X1 i_1807 (.ZN (n_2003), .A1 (inputB[9]), .A2 (inputA[28]));
INV_X1 i_1806 (.ZN (n_2002), .A (n_2003));
NAND3_X1 i_1805 (.ZN (n_2001), .A1 (inputB[8]), .A2 (inputA[27]), .A3 (n_2002));
NAND2_X1 i_1804 (.ZN (n_1999), .A1 (n_2004), .A2 (n_2001));
NAND2_X1 i_1803 (.ZN (n_1998), .A1 (inputB[10]), .A2 (inputA[26]));
XOR2_X1 i_1802 (.Z (n_4352), .A (n_1999), .B (n_1998));
NAND2_X1 i_1801 (.ZN (n_1997), .A1 (inputB[14]), .A2 (inputA[22]));
NOR2_X1 i_1800 (.ZN (n_1996), .A1 (n_2056), .A2 (n_1997));
AOI21_X1 i_1799 (.ZN (n_1995), .A (n_1996), .B1 (n_2056), .B2 (n_1997));
AND2_X1 i_1798 (.ZN (n_1992), .A1 (inputB[16]), .A2 (inputA[20]));
XOR2_X1 i_1797 (.Z (n_4338), .A (n_1995), .B (n_1992));
AOI22_X1 i_1795 (.ZN (n_1991), .A1 (inputB[18]), .A2 (inputA[18]), .B1 (inputB[17]), .B2 (inputA[19]));
INV_X1 i_1794 (.ZN (n_1990), .A (n_1991));
NAND4_X1 i_1793 (.ZN (n_1989), .A1 (inputB[18]), .A2 (inputA[18]), .A3 (inputB[17]), .A4 (inputA[19]));
NAND2_X1 i_1791 (.ZN (n_1988), .A1 (n_1990), .A2 (n_1989));
NAND2_X1 i_1790 (.ZN (n_1986), .A1 (inputB[19]), .A2 (inputA[17]));
XOR2_X1 i_1789 (.Z (n_4331), .A (n_1988), .B (n_1986));
NAND2_X1 i_1787 (.ZN (n_1985), .A1 (inputB[23]), .A2 (inputA[13]));
NOR2_X1 i_1786 (.ZN (n_1984), .A1 (n_2070), .A2 (n_1985));
AOI21_X1 i_1785 (.ZN (n_1980), .A (n_1984), .B1 (n_2070), .B2 (n_1985));
AND2_X1 i_1783 (.ZN (n_1975), .A1 (inputB[25]), .A2 (inputA[11]));
XOR2_X1 i_1782 (.Z (n_4317), .A (n_1980), .B (n_1975));
AOI22_X1 i_1781 (.ZN (n_1974), .A1 (inputB[27]), .A2 (inputA[9]), .B1 (inputB[26]), .B2 (inputA[10]));
INV_X1 i_1779 (.ZN (n_1970), .A (n_1974));
NAND3_X1 i_1778 (.ZN (n_1965), .A1 (inputB[27]), .A2 (inputA[10]), .A3 (n_2114));
NAND2_X1 i_1777 (.ZN (n_1964), .A1 (n_1970), .A2 (n_1965));
NAND2_X1 i_1775 (.ZN (n_1960), .A1 (inputB[28]), .A2 (inputA[8]));
XOR2_X1 i_1774 (.Z (n_4310), .A (n_1964), .B (n_1960));
AOI21_X1 i_1773 (.ZN (n_1955), .A (n_4226), .B1 (n_4225), .B2 (n_2080));
INV_X1 i_1771 (.ZN (n_4229), .A (n_1955));
NAND2_X1 i_1770 (.ZN (n_1954), .A1 (n_2105), .A2 (n_2103));
NAND2_X1 i_1769 (.ZN (n_1950), .A1 (n_2106), .A2 (n_1954));
XOR2_X1 i_1767 (.Z (n_4377), .A (n_4375), .B (n_1950));
OAI21_X1 i_1766 (.ZN (n_1945), .A (n_2132), .B1 (n_2135), .B2 (n_2130));
XOR2_X1 i_1765 (.Z (n_4367), .A (n_4365), .B (n_1945));
AOI21_X1 i_1763 (.ZN (n_1940), .A (n_4241), .B1 (n_4240), .B2 (n_2057));
INV_X1 i_1762 (.ZN (n_4244), .A (n_1940));
AOI21_X1 i_1761 (.ZN (n_1939), .A (n_4231), .B1 (n_4230), .B2 (n_2086));
INV_X1 i_1759 (.ZN (n_4234), .A (n_1939));
AOI21_X1 i_1758 (.ZN (n_1935), .A (n_4246), .B1 (n_4245), .B2 (n_2029));
INV_X1 i_1757 (.ZN (n_4249), .A (n_1935));
AOI21_X1 i_1756 (.ZN (n_1931), .A (n_4256), .B1 (n_4255), .B2 (n_2036));
INV_X1 i_1755 (.ZN (n_4259), .A (n_1931));
AOI21_X1 i_1754 (.ZN (n_1930), .A (n_4251), .B1 (n_4250), .B2 (n_2032));
INV_X1 i_1753 (.ZN (n_4254), .A (n_1930));
AND2_X1 i_1752 (.ZN (n_1929), .A1 (inputB[21]), .A2 (inputA[16]));
NAND2_X1 i_1751 (.ZN (n_1928), .A1 (n_2123), .A2 (n_1929));
AOI22_X1 i_1750 (.ZN (n_1927), .A1 (inputB[21]), .A2 (inputA[15]), .B1 (inputB[20]), .B2 (inputA[16]));
INV_X1 i_1749 (.ZN (n_1924), .A (n_1927));
NAND2_X1 i_1748 (.ZN (n_1923), .A1 (n_1928), .A2 (n_1924));
NAND2_X1 i_1747 (.ZN (n_1922), .A1 (inputB[22]), .A2 (inputA[14]));
XOR2_X1 i_1746 (.Z (n_1921), .A (n_1923), .B (n_1922));
XOR2_X1 i_1745 (.Z (n_4392), .A (n_4390), .B (n_1921));
NAND2_X1 i_1744 (.ZN (n_1919), .A1 (inputB[12]), .A2 (inputA[25]));
INV_X1 i_1743 (.ZN (n_1918), .A (n_1919));
NAND2_X1 i_1742 (.ZN (n_1917), .A1 (n_2136), .A2 (n_1918));
AOI22_X1 i_1741 (.ZN (n_1916), .A1 (inputB[12]), .A2 (inputA[24]), .B1 (inputB[11]), .B2 (inputA[25]));
INV_X1 i_1740 (.ZN (n_1915), .A (n_1916));
NAND2_X1 i_1739 (.ZN (n_1914), .A1 (n_1917), .A2 (n_1915));
NAND2_X1 i_1738 (.ZN (n_1911), .A1 (inputB[13]), .A2 (inputA[23]));
XOR2_X1 i_1737 (.Z (n_1910), .A (n_1914), .B (n_1911));
XOR2_X1 i_1736 (.Z (n_4387), .A (n_4385), .B (n_1910));
AOI21_X1 i_1735 (.ZN (n_1909), .A (n_4236), .B1 (n_4235), .B2 (n_2042));
INV_X1 i_1734 (.ZN (n_1908), .A (n_1909));
XNOR2_X1 i_1733 (.ZN (n_4407), .A (n_4405), .B (n_1909));
OAI21_X1 i_1732 (.ZN (n_1907), .A (n_2118), .B1 (n_2122), .B2 (n_2116));
XOR2_X1 i_1731 (.Z (n_1906), .A (n_4370), .B (n_1907));
XOR2_X1 i_1730 (.Z (n_4402), .A (n_4400), .B (n_1906));
AOI21_X1 i_1729 (.ZN (n_1904), .A (n_4211), .B1 (n_4210), .B2 (n_2035));
INV_X1 i_1728 (.ZN (n_1903), .A (n_1904));
XNOR2_X1 i_1727 (.ZN (n_1902), .A (n_4380), .B (n_1904));
XOR2_X1 i_1726 (.Z (n_4412), .A (n_4410), .B (n_1902));
AOI21_X1 i_1725 (.ZN (n_1901), .A (n_4271), .B1 (n_4270), .B2 (n_2025));
INV_X1 i_1724 (.ZN (n_4274), .A (n_1901));
AOI21_X1 i_1723 (.ZN (n_1900), .A (n_4276), .B1 (n_4275), .B2 (n_2023));
INV_X1 i_1722 (.ZN (n_4279), .A (n_1900));
AOI21_X1 i_1721 (.ZN (n_1898), .A (n_4102), .B1 (n_4101), .B2 (n_2210));
INV_X1 i_1720 (.ZN (n_1897), .A (n_1898));
AOI21_X1 i_1719 (.ZN (n_1896), .A (n_4261), .B1 (n_4260), .B2 (n_1897));
INV_X1 i_1718 (.ZN (n_1895), .A (n_1896));
XNOR2_X1 i_1717 (.ZN (n_4422), .A (n_4420), .B (n_1896));
AOI21_X1 i_1716 (.ZN (n_1894), .A (n_4266), .B1 (n_4265), .B2 (n_2028));
INV_X1 i_1715 (.ZN (n_1893), .A (n_1894));
XNOR2_X1 i_1714 (.ZN (n_4427), .A (n_4425), .B (n_1894));
NAND2_X1 i_1713 (.ZN (n_1890), .A1 (inputB[30]), .A2 (inputA[7]));
INV_X1 i_1712 (.ZN (n_1889), .A (n_1890));
AOI22_X1 i_1711 (.ZN (n_1888), .A1 (inputB[30]), .A2 (inputA[6]), .B1 (inputB[29]), .B2 (inputA[7]));
AOI21_X1 i_1710 (.ZN (n_1887), .A (n_1888), .B1 (n_2108), .B2 (n_1889));
NAND2_X1 i_1708 (.ZN (n_1886), .A1 (inputB[31]), .A2 (inputA[5]));
XOR2_X1 i_1707 (.Z (n_1885), .A (n_1887), .B (n_1886));
XOR2_X1 i_1706 (.Z (n_1883), .A (n_4395), .B (n_1885));
XOR2_X1 i_1704 (.Z (n_1882), .A (n_4415), .B (n_1883));
XOR2_X1 i_1703 (.Z (n_4432), .A (n_4430), .B (n_1882));
XNOR2_X1 i_1702 (.ZN (n_1878), .A (n_4260), .B (n_1898));
AOI21_X1 i_1700 (.ZN (n_1873), .A (n_4281), .B1 (n_4280), .B2 (n_1878));
INV_X1 i_1699 (.ZN (n_1872), .A (n_1873));
XNOR2_X1 i_1698 (.ZN (n_4437), .A (n_4435), .B (n_1873));
XOR2_X1 i_1696 (.Z (n_1868), .A (n_4280), .B (n_1878));
AOI21_X1 i_1695 (.ZN (n_1864), .A (n_4291), .B1 (n_4290), .B2 (n_1868));
INV_X1 i_1694 (.ZN (n_4294), .A (n_1864));
OAI21_X1 i_1692 (.ZN (n_4353), .A (n_2001), .B1 (n_2005), .B2 (n_1998));
OAI21_X1 i_1691 (.ZN (n_4346), .A (n_1917), .B1 (n_1916), .B2 (n_1911));
OAI21_X1 i_1690 (.ZN (n_4332), .A (n_1989), .B1 (n_1991), .B2 (n_1986));
OAI21_X1 i_1688 (.ZN (n_4325), .A (n_1928), .B1 (n_1927), .B2 (n_1922));
OAI21_X1 i_1687 (.ZN (n_4311), .A (n_1965), .B1 (n_1974), .B2 (n_1960));
AOI22_X1 i_1686 (.ZN (n_1863), .A1 (n_2108), .A2 (n_1889), .B1 (n_1887), .B2 (n_1886));
INV_X1 i_1684 (.ZN (n_4302), .A (n_1863));
AOI21_X1 i_1683 (.ZN (n_1862), .A (n_4371), .B1 (n_4370), .B2 (n_1907));
INV_X1 i_1682 (.ZN (n_4374), .A (n_1862));
AOI21_X1 i_1680 (.ZN (n_1858), .A (n_4366), .B1 (n_4365), .B2 (n_1945));
INV_X1 i_1679 (.ZN (n_4369), .A (n_1858));
NAND2_X1 i_1678 (.ZN (n_1853), .A1 (inputB[8]), .A2 (inputA[29]));
INV_X1 i_1676 (.ZN (n_1848), .A (n_1853));
NAND2_X1 i_1675 (.ZN (n_1847), .A1 (n_2002), .A2 (n_1848));
OAI21_X1 i_1674 (.ZN (n_1844), .A (n_1847), .B1 (n_2002), .B2 (n_1848));
NAND2_X1 i_1672 (.ZN (n_1843), .A1 (inputB[10]), .A2 (inputA[27]));
XOR2_X1 i_1671 (.Z (n_4502), .A (n_1844), .B (n_1843));
NAND2_X1 i_1670 (.ZN (n_1839), .A1 (inputB[11]), .A2 (inputA[26]));
INV_X1 i_1669 (.ZN (n_1838), .A (n_1839));
NAND2_X1 i_1668 (.ZN (n_1834), .A1 (n_1918), .A2 (n_1838));
OAI21_X1 i_1667 (.ZN (n_1833), .A (n_1834), .B1 (n_1918), .B2 (n_1838));
NAND2_X1 i_1666 (.ZN (n_1832), .A1 (inputB[13]), .A2 (inputA[24]));
XOR2_X1 i_1665 (.Z (n_4495), .A (n_1833), .B (n_1832));
AOI22_X1 i_1664 (.ZN (n_1831), .A1 (inputB[18]), .A2 (inputA[19]), .B1 (inputB[17]), .B2 (inputA[20]));
INV_X1 i_1663 (.ZN (n_1828), .A (n_1831));
NAND4_X1 i_1662 (.ZN (n_1827), .A1 (inputB[18]), .A2 (inputA[19]), .A3 (inputB[17]), .A4 (inputA[20]));
NAND2_X1 i_1661 (.ZN (n_1826), .A1 (n_1828), .A2 (n_1827));
NAND2_X1 i_1660 (.ZN (n_1825), .A1 (inputB[19]), .A2 (inputA[18]));
XOR2_X1 i_1659 (.Z (n_4481), .A (n_1826), .B (n_1825));
AOI21_X1 i_1658 (.ZN (n_1824), .A (n_1929), .B1 (inputB[20]), .B2 (inputA[17]));
INV_X1 i_1657 (.ZN (n_1823), .A (n_1824));
NAND3_X1 i_1656 (.ZN (n_1822), .A1 (inputB[20]), .A2 (inputA[17]), .A3 (n_1929));
NAND2_X1 i_1655 (.ZN (n_1821), .A1 (n_1823), .A2 (n_1822));
NAND2_X1 i_1654 (.ZN (n_1820), .A1 (inputB[22]), .A2 (inputA[15]));
XOR2_X1 i_1653 (.Z (n_4474), .A (n_1821), .B (n_1820));
AOI22_X1 i_1652 (.ZN (n_1819), .A1 (inputB[27]), .A2 (inputA[10]), .B1 (inputB[26]), .B2 (inputA[11]));
INV_X1 i_1651 (.ZN (n_1818), .A (n_1819));
NAND4_X1 i_1650 (.ZN (n_1817), .A1 (inputB[26]), .A2 (inputA[10]), .A3 (inputB[27]), .A4 (inputA[11]));
NAND2_X1 i_1649 (.ZN (n_1814), .A1 (n_1818), .A2 (n_1817));
NAND2_X1 i_1648 (.ZN (n_1813), .A1 (inputB[28]), .A2 (inputA[9]));
XOR2_X1 i_1647 (.Z (n_4460), .A (n_1814), .B (n_1813));
NAND2_X1 i_1646 (.ZN (n_1812), .A1 (inputB[29]), .A2 (inputA[8]));
INV_X1 i_1645 (.ZN (n_1811), .A (n_1812));
NAND2_X1 i_1644 (.ZN (n_1810), .A1 (n_1889), .A2 (n_1811));
NAND2_X1 i_1643 (.ZN (n_1807), .A1 (n_1890), .A2 (n_1812));
AND2_X1 i_1642 (.ZN (n_1806), .A1 (n_1810), .A2 (n_1807));
NAND2_X1 i_1641 (.ZN (n_1805), .A1 (inputB[31]), .A2 (inputA[6]));
XOR2_X1 i_1640 (.Z (n_4451), .A (n_1806), .B (n_1805));
AOI21_X1 i_1639 (.ZN (n_1804), .A (n_4376), .B1 (n_4375), .B2 (n_1950));
INV_X1 i_1638 (.ZN (n_1803), .A (n_1804));
XNOR2_X1 i_1637 (.ZN (n_4527), .A (n_4525), .B (n_1804));
NOR2_X1 i_1636 (.ZN (n_1802), .A1 (n_1984), .A2 (n_1975));
AOI21_X1 i_1635 (.ZN (n_1801), .A (n_1802), .B1 (n_2070), .B2 (n_1985));
XOR2_X1 i_1634 (.Z (n_4522), .A (n_4520), .B (n_1801));
AOI21_X1 i_1633 (.ZN (n_1800), .A (n_4396), .B1 (n_4395), .B2 (n_1885));
INV_X1 i_1632 (.ZN (n_4399), .A (n_1800));
AOI21_X1 i_1631 (.ZN (n_1799), .A (n_4391), .B1 (n_4390), .B2 (n_1921));
INV_X1 i_1629 (.ZN (n_4394), .A (n_1799));
AOI21_X1 i_1628 (.ZN (n_1798), .A (n_2009), .B1 (n_2010), .B2 (n_2006));
INV_X1 i_1627 (.ZN (n_1797), .A (n_1798));
NAND2_X1 i_1625 (.ZN (n_1796), .A1 (inputB[7]), .A2 (inputA[30]));
NAND2_X1 i_1624 (.ZN (n_1793), .A1 (inputB[6]), .A2 (inputA[31]));
XNOR2_X1 i_1623 (.ZN (n_1792), .A (n_1796), .B (n_1793));
XOR2_X1 i_1621 (.Z (n_1791), .A (n_1798), .B (n_1792));
XOR2_X1 i_1620 (.Z (n_4532), .A (n_4530), .B (n_1791));
AOI21_X1 i_1619 (.ZN (n_1790), .A (n_4406), .B1 (n_4405), .B2 (n_1908));
INV_X1 i_1617 (.ZN (n_4409), .A (n_1790));
AOI21_X1 i_1616 (.ZN (n_1789), .A (n_4381), .B1 (n_4380), .B2 (n_1903));
INV_X1 i_1615 (.ZN (n_1786), .A (n_1789));
XNOR2_X1 i_1613 (.ZN (n_4547), .A (n_4545), .B (n_1789));
AND2_X1 i_1612 (.ZN (n_1785), .A1 (inputB[24]), .A2 (inputA[14]));
NAND3_X1 i_1611 (.ZN (n_1781), .A1 (inputB[23]), .A2 (inputA[13]), .A3 (n_1785));
AOI22_X1 i_1609 (.ZN (n_1776), .A1 (inputB[24]), .A2 (inputA[13]), .B1 (inputB[23]), .B2 (inputA[14]));
INV_X1 i_1608 (.ZN (n_1775), .A (n_1776));
NAND2_X1 i_1607 (.ZN (n_1771), .A1 (n_1781), .A2 (n_1775));
NAND2_X1 i_1605 (.ZN (n_1767), .A1 (inputB[25]), .A2 (inputA[12]));
XOR2_X1 i_1604 (.Z (n_1766), .A (n_1771), .B (n_1767));
XOR2_X1 i_1603 (.Z (n_4542), .A (n_4540), .B (n_1766));
AOI21_X1 i_1601 (.ZN (n_1761), .A (n_4411), .B1 (n_4410), .B2 (n_1902));
INV_X1 i_1600 (.ZN (n_4414), .A (n_1761));
AOI21_X1 i_1599 (.ZN (n_1757), .A (n_4386), .B1 (n_4385), .B2 (n_1910));
INV_X1 i_1597 (.ZN (n_1756), .A (n_1757));
XNOR2_X1 i_1596 (.ZN (n_4557), .A (n_4555), .B (n_1757));
AOI21_X1 i_1595 (.ZN (n_1751), .A (n_4416), .B1 (n_4415), .B2 (n_1883));
INV_X1 i_1594 (.ZN (n_4419), .A (n_1751));
AOI21_X1 i_1593 (.ZN (n_1750), .A (n_4421), .B1 (n_4420), .B2 (n_1895));
INV_X1 i_1592 (.ZN (n_4424), .A (n_1750));
AOI21_X1 i_1591 (.ZN (n_1747), .A (n_4426), .B1 (n_4425), .B2 (n_1893));
INV_X1 i_1590 (.ZN (n_4429), .A (n_1747));
NAND2_X1 i_1589 (.ZN (n_1746), .A1 (inputB[16]), .A2 (inputA[21]));
AOI22_X1 i_1588 (.ZN (n_1745), .A1 (inputB[15]), .A2 (inputA[22]), .B1 (inputB[14]), .B2 (inputA[23]));
NAND4_X1 i_1587 (.ZN (n_1741), .A1 (inputB[14]), .A2 (inputA[22]), .A3 (inputB[15]), .A4 (inputA[23]));
INV_X1 i_1586 (.ZN (n_1737), .A (n_1741));
NOR2_X1 i_1585 (.ZN (n_1736), .A1 (n_1745), .A2 (n_1737));
XNOR2_X1 i_1584 (.ZN (n_1735), .A (n_1746), .B (n_1736));
XOR2_X1 i_1583 (.Z (n_1734), .A (n_4535), .B (n_1735));
XOR2_X1 i_1582 (.Z (n_4567), .A (n_4565), .B (n_1734));
NOR2_X1 i_1581 (.ZN (n_1732), .A1 (n_1996), .A2 (n_1992));
AOI21_X1 i_1580 (.ZN (n_1731), .A (n_1732), .B1 (n_2056), .B2 (n_1997));
XOR2_X1 i_1579 (.Z (n_1730), .A (n_4515), .B (n_1731));
XOR2_X1 i_1578 (.Z (n_1729), .A (n_4550), .B (n_1730));
XOR2_X1 i_1577 (.Z (n_4572), .A (n_4570), .B (n_1729));
AOI21_X1 i_1576 (.ZN (n_1728), .A (n_4401), .B1 (n_4400), .B2 (n_1906));
INV_X1 i_1575 (.ZN (n_1727), .A (n_1728));
XNOR2_X1 i_1574 (.ZN (n_1726), .A (n_4560), .B (n_1728));
XOR2_X1 i_1573 (.Z (n_4577), .A (n_4575), .B (n_1726));
AOI21_X1 i_1572 (.ZN (n_1725), .A (n_4286), .B1 (n_4285), .B2 (n_2019));
INV_X1 i_1571 (.ZN (n_1724), .A (n_1725));
AOI21_X1 i_1570 (.ZN (n_1723), .A (n_4441), .B1 (n_4440), .B2 (n_1724));
INV_X1 i_1569 (.ZN (n_4444), .A (n_1723));
AOI21_X1 i_1568 (.ZN (n_1722), .A (n_4431), .B1 (n_4430), .B2 (n_1882));
INV_X1 i_1567 (.ZN (n_1721), .A (n_1722));
XNOR2_X1 i_1566 (.ZN (n_4582), .A (n_4580), .B (n_1722));
NAND2_X1 i_1565 (.ZN (n_383), .A1 (inputB[7]), .A2 (inputA[31]));
AOI22_X1 i_1564 (.ZN (n_4503), .A1 (n_2003), .A2 (n_1853), .B1 (n_1847), .B2 (n_1843));
OAI21_X1 i_1563 (.ZN (n_4489), .A (n_1741), .B1 (n_1746), .B2 (n_1745));
OAI21_X1 i_1562 (.ZN (n_4482), .A (n_1827), .B1 (n_1831), .B2 (n_1825));
OAI21_X1 i_1561 (.ZN (n_4468), .A (n_1781), .B1 (n_1776), .B2 (n_1767));
OAI21_X1 i_1560 (.ZN (n_4461), .A (n_1817), .B1 (n_1819), .B2 (n_1813));
AOI21_X1 i_1559 (.ZN (n_1718), .A (n_4521), .B1 (n_4520), .B2 (n_1801));
INV_X1 i_1558 (.ZN (n_4524), .A (n_1718));
AOI21_X1 i_1557 (.ZN (n_1717), .A (n_4516), .B1 (n_4515), .B2 (n_1731));
INV_X1 i_1556 (.ZN (n_4519), .A (n_1717));
AOI22_X1 i_1555 (.ZN (n_1716), .A1 (inputB[9]), .A2 (inputA[29]), .B1 (inputB[8]), .B2 (inputA[30]));
INV_X1 i_1553 (.ZN (n_1715), .A (n_1716));
NAND2_X1 i_1552 (.ZN (n_1714), .A1 (inputB[9]), .A2 (inputA[30]));
OAI21_X1 i_1551 (.ZN (n_1711), .A (n_1715), .B1 (n_1853), .B2 (n_1714));
NAND2_X1 i_1549 (.ZN (n_1710), .A1 (inputB[10]), .A2 (inputA[28]));
XOR2_X1 i_1548 (.Z (n_4647), .A (n_1711), .B (n_1710));
AOI22_X1 i_1547 (.ZN (n_1709), .A1 (inputB[12]), .A2 (inputA[26]), .B1 (inputB[11]), .B2 (inputA[27]));
INV_X1 i_1545 (.ZN (n_1708), .A (n_1709));
AND2_X1 i_1544 (.ZN (n_1707), .A1 (inputB[12]), .A2 (inputA[27]));
NAND2_X1 i_1543 (.ZN (n_1706), .A1 (n_1838), .A2 (n_1707));
NAND2_X1 i_1541 (.ZN (n_1705), .A1 (n_1708), .A2 (n_1706));
NAND2_X1 i_1540 (.ZN (n_1704), .A1 (inputB[13]), .A2 (inputA[25]));
XOR2_X1 i_1539 (.Z (n_4640), .A (n_1705), .B (n_1704));
AND2_X1 i_1537 (.ZN (n_1703), .A1 (inputB[17]), .A2 (inputA[21]));
AOI21_X1 i_1536 (.ZN (n_1702), .A (n_1703), .B1 (inputB[18]), .B2 (inputA[20]));
INV_X1 i_1535 (.ZN (n_1701), .A (n_1702));
NAND3_X1 i_1533 (.ZN (n_1700), .A1 (inputB[18]), .A2 (inputA[20]), .A3 (n_1703));
NAND2_X1 i_1532 (.ZN (n_1697), .A1 (n_1701), .A2 (n_1700));
NAND2_X1 i_1531 (.ZN (n_1696), .A1 (inputB[19]), .A2 (inputA[19]));
XOR2_X1 i_1529 (.Z (n_4626), .A (n_1697), .B (n_1696));
AND2_X1 i_1528 (.ZN (n_1692), .A1 (inputB[20]), .A2 (inputA[18]));
AOI21_X1 i_1527 (.ZN (n_1687), .A (n_1692), .B1 (inputB[21]), .B2 (inputA[17]));
INV_X1 i_1525 (.ZN (n_1686), .A (n_1687));
NAND3_X1 i_1524 (.ZN (n_1683), .A1 (inputB[21]), .A2 (inputA[17]), .A3 (n_1692));
NAND2_X1 i_1523 (.ZN (n_1682), .A1 (n_1686), .A2 (n_1683));
NAND2_X1 i_1522 (.ZN (n_1677), .A1 (inputB[22]), .A2 (inputA[16]));
XOR2_X1 i_1521 (.Z (n_4619), .A (n_1682), .B (n_1677));
AOI22_X1 i_1520 (.ZN (n_1672), .A1 (inputB[27]), .A2 (inputA[11]), .B1 (inputB[26]), .B2 (inputA[12]));
INV_X1 i_1519 (.ZN (n_1671), .A (n_1672));
NAND4_X1 i_1518 (.ZN (n_1668), .A1 (inputB[26]), .A2 (inputA[11]), .A3 (inputB[27]), .A4 (inputA[12]));
NAND2_X1 i_1517 (.ZN (n_1667), .A1 (n_1671), .A2 (n_1668));
NAND2_X1 i_1516 (.ZN (n_1662), .A1 (inputB[28]), .A2 (inputA[10]));
XOR2_X1 i_1515 (.Z (n_4605), .A (n_1667), .B (n_1662));
NAND2_X1 i_1514 (.ZN (n_1658), .A1 (inputB[30]), .A2 (inputA[9]));
INV_X1 i_1513 (.ZN (n_1657), .A (n_1658));
AOI22_X1 i_1512 (.ZN (n_1653), .A1 (inputB[30]), .A2 (inputA[8]), .B1 (inputB[29]), .B2 (inputA[9]));
AOI21_X1 i_1511 (.ZN (n_1652), .A (n_1653), .B1 (n_1811), .B2 (n_1657));
NAND2_X1 i_1510 (.ZN (n_1651), .A1 (inputB[31]), .A2 (inputA[7]));
XOR2_X1 i_1509 (.Z (n_4596), .A (n_1652), .B (n_1651));
NAND2_X1 i_1508 (.ZN (n_1650), .A1 (n_1807), .A2 (n_1805));
NAND2_X1 i_1507 (.ZN (n_1649), .A1 (n_1810), .A2 (n_1650));
XOR2_X1 i_1506 (.Z (n_4664), .A (n_4662), .B (n_1649));
OAI21_X1 i_1505 (.ZN (n_1646), .A (n_1822), .B1 (n_1824), .B2 (n_1820));
XOR2_X1 i_1504 (.Z (n_4659), .A (n_4657), .B (n_1646));
AOI21_X1 i_1503 (.ZN (n_1645), .A (n_4541), .B1 (n_4540), .B2 (n_1766));
INV_X1 i_1502 (.ZN (n_4544), .A (n_1645));
AOI21_X1 i_1501 (.ZN (n_1644), .A (n_4536), .B1 (n_4535), .B2 (n_1735));
INV_X1 i_1500 (.ZN (n_4539), .A (n_1644));
AOI21_X1 i_1499 (.ZN (n_1643), .A (n_4546), .B1 (n_4545), .B2 (n_1786));
INV_X1 i_1498 (.ZN (n_4549), .A (n_1643));
AOI21_X1 i_1497 (.ZN (n_1640), .A (n_1796), .B1 (n_1797), .B2 (n_1792));
AOI21_X1 i_1496 (.ZN (n_1639), .A (n_1640), .B1 (n_1798), .B2 (n_1793));
INV_X1 i_1495 (.ZN (n_1638), .A (n_1639));
XNOR2_X1 i_1494 (.ZN (n_4669), .A (n_4667), .B (n_1639));
AOI21_X1 i_1493 (.ZN (n_1637), .A (n_4551), .B1 (n_4550), .B2 (n_1730));
INV_X1 i_1492 (.ZN (n_4554), .A (n_1637));
AOI21_X1 i_1491 (.ZN (n_1636), .A (n_4526), .B1 (n_4525), .B2 (n_1803));
INV_X1 i_1490 (.ZN (n_1634), .A (n_1636));
XNOR2_X1 i_1489 (.ZN (n_4684), .A (n_4682), .B (n_1636));
AOI22_X1 i_1488 (.ZN (n_1633), .A1 (inputB[15]), .A2 (inputA[23]), .B1 (inputB[14]), .B2 (inputA[24]));
INV_X1 i_1487 (.ZN (n_1632), .A (n_1633));
NAND2_X1 i_1486 (.ZN (n_1631), .A1 (inputB[15]), .A2 (inputA[24]));
INV_X1 i_1485 (.ZN (n_1630), .A (n_1631));
NAND3_X1 i_1484 (.ZN (n_1629), .A1 (inputB[14]), .A2 (inputA[23]), .A3 (n_1630));
NAND2_X1 i_1483 (.ZN (n_1628), .A1 (n_1632), .A2 (n_1629));
NAND2_X1 i_1481 (.ZN (n_1626), .A1 (inputB[16]), .A2 (inputA[22]));
XOR2_X1 i_1480 (.Z (n_1625), .A (n_1628), .B (n_1626));
XOR2_X1 i_1479 (.Z (n_4674), .A (n_4672), .B (n_1625));
AOI21_X1 i_1477 (.ZN (n_1624), .A (n_4561), .B1 (n_4560), .B2 (n_1727));
INV_X1 i_1476 (.ZN (n_4564), .A (n_1624));
AOI22_X1 i_1475 (.ZN (n_1623), .A1 (n_1919), .A2 (n_1839), .B1 (n_1834), .B2 (n_1832));
XOR2_X1 i_1473 (.Z (n_1622), .A (n_4652), .B (n_1623));
XOR2_X1 i_1472 (.Z (n_4689), .A (n_4687), .B (n_1622));
AOI21_X1 i_1471 (.ZN (n_1619), .A (n_4566), .B1 (n_4565), .B2 (n_1734));
INV_X1 i_1469 (.ZN (n_4569), .A (n_1619));
AOI21_X1 i_1468 (.ZN (n_1618), .A (n_4571), .B1 (n_4570), .B2 (n_1729));
INV_X1 i_1467 (.ZN (n_4574), .A (n_1618));
AOI21_X1 i_1465 (.ZN (n_1617), .A (n_1785), .B1 (inputB[23]), .B2 (inputA[15]));
INV_X1 i_1464 (.ZN (n_1616), .A (n_1617));
NAND3_X1 i_1463 (.ZN (n_1615), .A1 (inputB[23]), .A2 (inputA[15]), .A3 (n_1785));
NAND2_X1 i_1461 (.ZN (n_1613), .A1 (n_1616), .A2 (n_1615));
NAND2_X1 i_1460 (.ZN (n_1612), .A1 (inputB[25]), .A2 (inputA[13]));
XOR2_X1 i_1459 (.Z (n_1611), .A (n_1613), .B (n_1612));
XOR2_X1 i_1457 (.Z (n_1607), .A (n_4677), .B (n_1611));
XOR2_X1 i_1456 (.Z (n_4704), .A (n_4702), .B (n_1607));
AOI21_X1 i_1455 (.ZN (n_1602), .A (n_4576), .B1 (n_4575), .B2 (n_1726));
INV_X1 i_1453 (.ZN (n_4579), .A (n_1602));
AOI21_X1 i_1452 (.ZN (n_1601), .A (n_4556), .B1 (n_4555), .B2 (n_1756));
INV_X1 i_1451 (.ZN (n_1598), .A (n_1601));
XNOR2_X1 i_1450 (.ZN (n_1597), .A (n_4697), .B (n_1601));
XOR2_X1 i_1449 (.Z (n_4714), .A (n_4712), .B (n_1597));
AOI21_X1 i_1448 (.ZN (n_1592), .A (n_4436), .B1 (n_4435), .B2 (n_1872));
INV_X1 i_1447 (.ZN (n_1591), .A (n_1592));
AOI21_X1 i_1446 (.ZN (n_1587), .A (n_4586), .B1 (n_4585), .B2 (n_1591));
INV_X1 i_1445 (.ZN (n_4589), .A (n_1587));
AOI21_X1 i_1444 (.ZN (n_1586), .A (n_4531), .B1 (n_4530), .B2 (n_1791));
INV_X1 i_1443 (.ZN (n_1583), .A (n_1586));
XNOR2_X1 i_1442 (.ZN (n_1582), .A (n_4692), .B (n_1586));
XOR2_X1 i_1441 (.Z (n_1577), .A (n_4707), .B (n_1582));
XOR2_X1 i_1440 (.Z (n_4719), .A (n_4717), .B (n_1577));
OAI22_X1 i_1439 (.ZN (n_4648), .A1 (n_1853), .A2 (n_1714), .B1 (n_1716), .B2 (n_1710));
OAI21_X1 i_1438 (.ZN (n_4641), .A (n_1706), .B1 (n_1709), .B2 (n_1704));
OAI21_X1 i_1437 (.ZN (n_4627), .A (n_1700), .B1 (n_1702), .B2 (n_1696));
OAI21_X1 i_1436 (.ZN (n_4620), .A (n_1683), .B1 (n_1687), .B2 (n_1677));
OAI21_X1 i_1435 (.ZN (n_4606), .A (n_1668), .B1 (n_1672), .B2 (n_1662));
AOI21_X1 i_1434 (.ZN (n_1573), .A (n_1651), .B1 (n_1811), .B2 (n_1657));
NOR2_X1 i_1433 (.ZN (n_4597), .A1 (n_1653), .A2 (n_1573));
AOI21_X1 i_1432 (.ZN (n_1572), .A (n_4658), .B1 (n_4657), .B2 (n_1646));
INV_X1 i_1431 (.ZN (n_4661), .A (n_1572));
AOI21_X1 i_1430 (.ZN (n_1571), .A (n_4653), .B1 (n_4652), .B2 (n_1623));
INV_X1 i_1429 (.ZN (n_4656), .A (n_1571));
AOI21_X1 i_1428 (.ZN (n_1570), .A (n_1707), .B1 (inputB[11]), .B2 (inputA[28]));
INV_X1 i_1427 (.ZN (n_1569), .A (n_1570));
NAND3_X1 i_1426 (.ZN (n_1568), .A1 (inputB[11]), .A2 (inputA[28]), .A3 (n_1707));
NAND2_X1 i_1425 (.ZN (n_1567), .A1 (n_1569), .A2 (n_1568));
NAND2_X1 i_1424 (.ZN (n_1566), .A1 (inputB[13]), .A2 (inputA[26]));
XOR2_X1 i_1423 (.Z (n_4777), .A (n_1567), .B (n_1566));
NAND2_X1 i_1422 (.ZN (n_1565), .A1 (inputB[14]), .A2 (inputA[25]));
INV_X1 i_1421 (.ZN (n_1564), .A (n_1565));
NAND2_X1 i_1420 (.ZN (n_1563), .A1 (n_1630), .A2 (n_1564));
OAI21_X1 i_1419 (.ZN (n_1562), .A (n_1563), .B1 (n_1630), .B2 (n_1564));
NAND2_X1 i_1417 (.ZN (n_1560), .A1 (inputB[16]), .A2 (inputA[23]));
XOR2_X1 i_1416 (.Z (n_4770), .A (n_1562), .B (n_1560));
AOI22_X1 i_1415 (.ZN (n_1559), .A1 (inputB[21]), .A2 (inputA[18]), .B1 (inputB[20]), .B2 (inputA[19]));
INV_X1 i_1413 (.ZN (n_1558), .A (n_1559));
NAND2_X1 i_1412 (.ZN (n_1557), .A1 (inputB[21]), .A2 (inputA[19]));
INV_X1 i_1411 (.ZN (n_1556), .A (n_1557));
NAND2_X1 i_1409 (.ZN (n_1554), .A1 (n_1692), .A2 (n_1556));
NAND2_X1 i_1408 (.ZN (n_1553), .A1 (n_1558), .A2 (n_1554));
NAND2_X1 i_1407 (.ZN (n_1552), .A1 (inputB[22]), .A2 (inputA[17]));
XOR2_X1 i_1405 (.Z (n_4756), .A (n_1553), .B (n_1552));
AND2_X1 i_1404 (.ZN (n_1551), .A1 (inputB[23]), .A2 (inputA[16]));
AOI21_X1 i_1403 (.ZN (n_1550), .A (n_1551), .B1 (inputB[24]), .B2 (inputA[15]));
INV_X1 i_1401 (.ZN (n_1549), .A (n_1550));
NAND3_X1 i_1400 (.ZN (n_1546), .A1 (inputB[24]), .A2 (inputA[15]), .A3 (n_1551));
NAND2_X1 i_1399 (.ZN (n_1545), .A1 (n_1549), .A2 (n_1546));
NAND2_X1 i_1397 (.ZN (n_1544), .A1 (inputB[25]), .A2 (inputA[14]));
XOR2_X1 i_1396 (.Z (n_4749), .A (n_1545), .B (n_1544));
NAND2_X1 i_1395 (.ZN (n_1543), .A1 (inputB[29]), .A2 (inputA[10]));
INV_X1 i_1393 (.ZN (n_1542), .A (n_1543));
NAND2_X1 i_1392 (.ZN (n_1541), .A1 (n_1657), .A2 (n_1542));
NAND2_X1 i_1391 (.ZN (n_1539), .A1 (n_1658), .A2 (n_1543));
AND2_X1 i_1390 (.ZN (n_1538), .A1 (n_1541), .A2 (n_1539));
NAND2_X1 i_1389 (.ZN (n_1537), .A1 (inputB[31]), .A2 (inputA[8]));
XOR2_X1 i_1388 (.Z (n_4733), .A (n_1538), .B (n_1537));
AOI21_X1 i_1387 (.ZN (n_1536), .A (n_4668), .B1 (n_4667), .B2 (n_1638));
INV_X1 i_1386 (.ZN (n_4671), .A (n_1536));
OAI21_X1 i_1385 (.ZN (n_1535), .A (n_1615), .B1 (n_1617), .B2 (n_1612));
XOR2_X1 i_1384 (.Z (n_4797), .A (n_4795), .B (n_1535));
OAI21_X1 i_1383 (.ZN (n_1533), .A (n_1629), .B1 (n_1633), .B2 (n_1626));
XOR2_X1 i_1382 (.Z (n_4792), .A (n_4790), .B (n_1533));
AOI21_X1 i_1381 (.ZN (n_1532), .A (n_4673), .B1 (n_4672), .B2 (n_1625));
INV_X1 i_1380 (.ZN (n_4676), .A (n_1532));
AOI21_X1 i_1379 (.ZN (n_1531), .A (n_4683), .B1 (n_4682), .B2 (n_1634));
INV_X1 i_1378 (.ZN (n_4686), .A (n_1531));
AOI21_X1 i_1377 (.ZN (n_1527), .A (n_4693), .B1 (n_4692), .B2 (n_1583));
INV_X1 i_1376 (.ZN (n_4696), .A (n_1527));
AOI21_X1 i_1375 (.ZN (n_1522), .A (n_4688), .B1 (n_4687), .B2 (n_1622));
INV_X1 i_1374 (.ZN (n_4691), .A (n_1522));
AND2_X1 i_1373 (.ZN (n_1521), .A1 (inputB[18]), .A2 (inputA[22]));
NAND2_X1 i_1372 (.ZN (n_1517), .A1 (n_1703), .A2 (n_1521));
AOI22_X1 i_1371 (.ZN (n_1512), .A1 (inputB[18]), .A2 (inputA[21]), .B1 (inputB[17]), .B2 (inputA[22]));
INV_X1 i_1370 (.ZN (n_1507), .A (n_1512));
NAND2_X1 i_1369 (.ZN (n_1506), .A1 (n_1517), .A2 (n_1507));
NAND2_X1 i_1368 (.ZN (n_1502), .A1 (inputB[19]), .A2 (inputA[20]));
XOR2_X1 i_1367 (.Z (n_1501), .A (n_1506), .B (n_1502));
XOR2_X1 i_1366 (.Z (n_4812), .A (n_4810), .B (n_1501));
AOI21_X1 i_1365 (.ZN (n_1497), .A (n_4663), .B1 (n_4662), .B2 (n_1649));
INV_X1 i_1364 (.ZN (n_1496), .A (n_1497));
XNOR2_X1 i_1363 (.ZN (n_1493), .A (n_4800), .B (n_1497));
XOR2_X1 i_1362 (.Z (n_4822), .A (n_4820), .B (n_1493));
AOI21_X1 i_1361 (.ZN (n_1492), .A (n_4678), .B1 (n_4677), .B2 (n_1611));
INV_X1 i_1360 (.ZN (n_1491), .A (n_1492));
XNOR2_X1 i_1359 (.ZN (n_4827), .A (n_4825), .B (n_1492));
AOI21_X1 i_1358 (.ZN (n_1490), .A (n_4703), .B1 (n_4702), .B2 (n_1607));
INV_X1 i_1356 (.ZN (n_4706), .A (n_1490));
AOI22_X1 i_1355 (.ZN (n_1488), .A1 (inputB[27]), .A2 (inputA[12]), .B1 (inputB[26]), .B2 (inputA[13]));
INV_X1 i_1354 (.ZN (n_1487), .A (n_1488));
NAND4_X1 i_1352 (.ZN (n_1486), .A1 (inputB[26]), .A2 (inputA[12]), .A3 (inputB[27]), .A4 (inputA[13]));
NAND2_X1 i_1351 (.ZN (n_1485), .A1 (n_1487), .A2 (n_1486));
NAND2_X1 i_1350 (.ZN (n_1484), .A1 (inputB[28]), .A2 (inputA[11]));
XOR2_X1 i_1348 (.Z (n_1483), .A (n_1485), .B (n_1484));
XOR2_X1 i_1347 (.Z (n_1481), .A (n_4815), .B (n_1483));
XOR2_X1 i_1346 (.Z (n_4837), .A (n_4835), .B (n_1481));
AOI21_X1 i_1344 (.ZN (n_1480), .A (n_4708), .B1 (n_4707), .B2 (n_1582));
INV_X1 i_1343 (.ZN (n_4711), .A (n_1480));
AOI21_X1 i_1342 (.ZN (n_1479), .A (n_4713), .B1 (n_4712), .B2 (n_1597));
INV_X1 i_1340 (.ZN (n_4716), .A (n_1479));
AND3_X1 i_1339 (.ZN (n_1478), .A1 (inputB[8]), .A2 (inputA[31]), .A3 (n_1714));
AOI21_X1 i_1338 (.ZN (n_1477), .A (n_1714), .B1 (inputB[8]), .B2 (inputA[31]));
INV_X1 i_1336 (.ZN (n_1475), .A (n_1477));
NOR2_X1 i_1335 (.ZN (n_1474), .A1 (n_1478), .A2 (n_1477));
NAND2_X1 i_1334 (.ZN (n_1473), .A1 (inputB[10]), .A2 (inputA[29]));
XNOR2_X1 i_1333 (.ZN (n_1472), .A (n_1474), .B (n_1473));
XOR2_X1 i_1332 (.Z (n_1471), .A (n_4805), .B (n_1472));
XOR2_X1 i_1331 (.Z (n_1470), .A (n_4830), .B (n_1471));
XOR2_X1 i_1330 (.Z (n_4847), .A (n_4845), .B (n_1470));
AOI21_X1 i_1329 (.ZN (n_1467), .A (n_4698), .B1 (n_4697), .B2 (n_1598));
INV_X1 i_1328 (.ZN (n_1466), .A (n_1467));
XNOR2_X1 i_1327 (.ZN (n_1465), .A (n_4840), .B (n_1467));
XOR2_X1 i_1326 (.Z (n_4852), .A (n_4850), .B (n_1465));
AOI21_X1 i_1325 (.ZN (n_1464), .A (n_4581), .B1 (n_4580), .B2 (n_1721));
INV_X1 i_1324 (.ZN (n_1463), .A (n_1464));
AOI21_X1 i_1323 (.ZN (n_1462), .A (n_4723), .B1 (n_4722), .B2 (n_1463));
INV_X1 i_1322 (.ZN (n_4726), .A (n_1462));
OAI21_X1 i_1321 (.ZN (n_4778), .A (n_1568), .B1 (n_1570), .B2 (n_1566));
AOI22_X1 i_1320 (.ZN (n_4771), .A1 (n_1631), .A2 (n_1565), .B1 (n_1563), .B2 (n_1560));
OAI21_X1 i_1319 (.ZN (n_4757), .A (n_1554), .B1 (n_1559), .B2 (n_1552));
OAI21_X1 i_1318 (.ZN (n_4750), .A (n_1546), .B1 (n_1550), .B2 (n_1544));
NAND2_X1 i_1317 (.ZN (n_1460), .A1 (n_1539), .A2 (n_1537));
NAND2_X1 i_1316 (.ZN (n_4734), .A1 (n_1541), .A2 (n_1460));
AOI21_X1 i_1315 (.ZN (n_1459), .A (n_4796), .B1 (n_4795), .B2 (n_1535));
INV_X1 i_1314 (.ZN (n_4799), .A (n_1459));
AOI211_X1 i_1313 (.ZN (n_1455), .A (n_5757), .B (n_5753), .C1 (inputB[10]), .C2 (inputA[30]));
OAI211_X1 i_1312 (.ZN (n_1450), .A (inputB[10]), .B (inputA[30]), .C1 (n_5757), .C2 (n_5753));
INV_X1 i_1311 (.ZN (n_1445), .A (n_1450));
NOR2_X1 i_1310 (.ZN (n_1440), .A1 (n_1455), .A2 (n_1445));
AOI21_X1 i_1309 (.ZN (n_1435), .A (n_1478), .B1 (n_1475), .B2 (n_1473));
INV_X1 i_1308 (.ZN (n_1434), .A (n_1435));
XOR2_X1 i_1307 (.Z (n_4917), .A (n_1440), .B (n_1435));
NOR2_X1 i_1306 (.ZN (n_1430), .A1 (n_5758), .A2 (n_5750));
AOI21_X1 i_1305 (.ZN (n_1426), .A (n_1430), .B1 (inputB[12]), .B2 (inputA[28]));
INV_X1 i_1304 (.ZN (n_1425), .A (n_1426));
NAND3_X1 i_1303 (.ZN (n_1424), .A1 (inputB[12]), .A2 (inputA[28]), .A3 (n_1430));
NAND2_X1 i_1302 (.ZN (n_1423), .A1 (n_1425), .A2 (n_1424));
NAND2_X1 i_1301 (.ZN (n_1422), .A1 (inputB[13]), .A2 (inputA[27]));
XOR2_X1 i_1299 (.Z (n_4910), .A (n_1423), .B (n_1422));
AOI21_X1 i_1298 (.ZN (n_1421), .A (n_1521), .B1 (inputB[17]), .B2 (inputA[23]));
INV_X1 i_1297 (.ZN (n_1419), .A (n_1421));
NAND3_X1 i_1295 (.ZN (n_1418), .A1 (inputB[17]), .A2 (inputA[23]), .A3 (n_1521));
NAND2_X1 i_1294 (.ZN (n_1417), .A1 (n_1419), .A2 (n_1418));
NAND2_X1 i_1293 (.ZN (n_1416), .A1 (inputB[19]), .A2 (inputA[21]));
XOR2_X1 i_1291 (.Z (n_4896), .A (n_1417), .B (n_1416));
NAND2_X1 i_1290 (.ZN (n_1414), .A1 (inputB[20]), .A2 (inputA[20]));
INV_X1 i_1289 (.ZN (n_1413), .A (n_1414));
NAND2_X1 i_1287 (.ZN (n_1412), .A1 (n_1556), .A2 (n_1413));
OAI21_X1 i_1286 (.ZN (n_1411), .A (n_1412), .B1 (n_1556), .B2 (n_1413));
NAND2_X1 i_1285 (.ZN (n_1410), .A1 (inputB[22]), .A2 (inputA[18]));
XOR2_X1 i_1283 (.Z (n_4889), .A (n_1411), .B (n_1410));
AOI22_X1 i_1282 (.ZN (n_1409), .A1 (inputB[27]), .A2 (inputA[13]), .B1 (inputB[26]), .B2 (inputA[14]));
INV_X1 i_1281 (.ZN (n_1406), .A (n_1409));
NAND2_X1 i_1279 (.ZN (n_1405), .A1 (inputB[27]), .A2 (inputA[14]));
INV_X1 i_1278 (.ZN (n_1404), .A (n_1405));
NAND3_X1 i_1277 (.ZN (n_1403), .A1 (inputB[26]), .A2 (inputA[13]), .A3 (n_1404));
NAND2_X1 i_1276 (.ZN (n_1402), .A1 (n_1406), .A2 (n_1403));
NAND2_X1 i_1275 (.ZN (n_1401), .A1 (inputB[28]), .A2 (inputA[12]));
XOR2_X1 i_1274 (.Z (n_4875), .A (n_1402), .B (n_1401));
AOI22_X1 i_1273 (.ZN (n_1399), .A1 (inputB[30]), .A2 (inputA[10]), .B1 (inputB[29]), .B2 (inputA[11]));
INV_X1 i_1272 (.ZN (n_1398), .A (n_1399));
NAND3_X1 i_1271 (.ZN (n_1397), .A1 (inputB[30]), .A2 (inputA[11]), .A3 (n_1542));
NAND2_X1 i_1270 (.ZN (n_1396), .A1 (n_1398), .A2 (n_1397));
AND2_X1 i_1269 (.ZN (n_1395), .A1 (inputB[31]), .A2 (inputA[9]));
XOR2_X1 i_1268 (.Z (n_4866), .A (n_1396), .B (n_1395));
OAI21_X1 i_1267 (.ZN (n_1393), .A (n_1486), .B1 (n_1488), .B2 (n_1484));
XOR2_X1 i_1266 (.Z (n_4930), .A (n_4928), .B (n_1393));
AOI21_X1 i_1265 (.ZN (n_1392), .A (n_1512), .B1 (n_1517), .B2 (n_1502));
XOR2_X1 i_1264 (.Z (n_4925), .A (n_4923), .B (n_1392));
AOI21_X1 i_1263 (.ZN (n_1391), .A (n_4811), .B1 (n_4810), .B2 (n_1501));
INV_X1 i_1262 (.ZN (n_4814), .A (n_1391));
AOI21_X1 i_1261 (.ZN (n_1388), .A (n_4806), .B1 (n_4805), .B2 (n_1472));
INV_X1 i_1260 (.ZN (n_4809), .A (n_1388));
AOI21_X1 i_1259 (.ZN (n_1387), .A (n_4826), .B1 (n_4825), .B2 (n_1491));
INV_X1 i_1258 (.ZN (n_4829), .A (n_1387));
AOI21_X1 i_1257 (.ZN (n_1382), .A (n_4821), .B1 (n_4820), .B2 (n_1493));
INV_X1 i_1256 (.ZN (n_4824), .A (n_1382));
NAND3_X1 i_1255 (.ZN (n_1381), .A1 (inputB[24]), .A2 (inputA[17]), .A3 (n_1551));
AOI22_X1 i_1254 (.ZN (n_1377), .A1 (inputB[24]), .A2 (inputA[16]), .B1 (inputB[23]), .B2 (inputA[17]));
INV_X1 i_1253 (.ZN (n_1373), .A (n_1377));
NAND2_X1 i_1252 (.ZN (n_1372), .A1 (n_1381), .A2 (n_1373));
NAND2_X1 i_1250 (.ZN (n_1371), .A1 (inputB[25]), .A2 (inputA[15]));
XOR2_X1 i_1249 (.Z (n_1367), .A (n_1372), .B (n_1371));
XOR2_X1 i_1248 (.Z (n_4945), .A (n_4943), .B (n_1367));
AOI22_X1 i_1246 (.ZN (n_1363), .A1 (inputB[15]), .A2 (inputA[25]), .B1 (inputB[14]), .B2 (inputA[26]));
INV_X1 i_1245 (.ZN (n_1362), .A (n_1363));
AND2_X1 i_1244 (.ZN (n_1361), .A1 (inputB[15]), .A2 (inputA[26]));
NAND2_X1 i_1242 (.ZN (n_1360), .A1 (n_1564), .A2 (n_1361));
NAND2_X1 i_1241 (.ZN (n_1358), .A1 (n_1362), .A2 (n_1360));
NAND2_X1 i_1240 (.ZN (n_1357), .A1 (inputB[16]), .A2 (inputA[24]));
XOR2_X1 i_1238 (.Z (n_1356), .A (n_1358), .B (n_1357));
XOR2_X1 i_1237 (.Z (n_4940), .A (n_4938), .B (n_1356));
AOI21_X1 i_1236 (.ZN (n_1355), .A (n_4791), .B1 (n_4790), .B2 (n_1533));
INV_X1 i_1234 (.ZN (n_1354), .A (n_1355));
XNOR2_X1 i_1233 (.ZN (n_1353), .A (n_4933), .B (n_1355));
XOR2_X1 i_1232 (.Z (n_4960), .A (n_4958), .B (n_1353));
AOI21_X1 i_1231 (.ZN (n_1352), .A (n_4816), .B1 (n_4815), .B2 (n_1483));
INV_X1 i_1230 (.ZN (n_1350), .A (n_1352));
XNOR2_X1 i_1229 (.ZN (n_4955), .A (n_4953), .B (n_1352));
AOI21_X1 i_1228 (.ZN (n_1349), .A (n_4841), .B1 (n_4840), .B2 (n_1466));
INV_X1 i_1227 (.ZN (n_4844), .A (n_1349));
AOI21_X1 i_1226 (.ZN (n_1348), .A (n_4801), .B1 (n_4800), .B2 (n_1496));
INV_X1 i_1225 (.ZN (n_1347), .A (n_1348));
XNOR2_X1 i_1224 (.ZN (n_1346), .A (n_4948), .B (n_1348));
XOR2_X1 i_1223 (.Z (n_4965), .A (n_4963), .B (n_1346));
AOI21_X1 i_1222 (.ZN (n_1343), .A (n_4831), .B1 (n_4830), .B2 (n_1471));
INV_X1 i_1221 (.ZN (n_1342), .A (n_1343));
XNOR2_X1 i_1220 (.ZN (n_4970), .A (n_4968), .B (n_1343));
AOI21_X1 i_1219 (.ZN (n_1341), .A (n_4836), .B1 (n_4835), .B2 (n_1481));
INV_X1 i_1218 (.ZN (n_1340), .A (n_1341));
XNOR2_X1 i_1217 (.ZN (n_4975), .A (n_4973), .B (n_1341));
AOI21_X1 i_1216 (.ZN (n_1339), .A (n_4846), .B1 (n_4845), .B2 (n_1470));
INV_X1 i_1215 (.ZN (n_1337), .A (n_1339));
XNOR2_X1 i_1214 (.ZN (n_4980), .A (n_4978), .B (n_1339));
AOI21_X1 i_1213 (.ZN (n_1336), .A (n_4718), .B1 (n_4717), .B2 (n_1577));
INV_X1 i_1212 (.ZN (n_1335), .A (n_1336));
AOI21_X1 i_1211 (.ZN (n_1334), .A (n_4856), .B1 (n_4855), .B2 (n_1335));
INV_X1 i_1210 (.ZN (n_4859), .A (n_1334));
NAND2_X1 i_1209 (.ZN (n_382), .A1 (inputB[10]), .A2 (inputA[31]));
OAI21_X1 i_1208 (.ZN (n_4911), .A (n_1424), .B1 (n_1426), .B2 (n_1422));
OAI21_X1 i_1207 (.ZN (n_4897), .A (n_1418), .B1 (n_1421), .B2 (n_1416));
AOI22_X1 i_1206 (.ZN (n_4890), .A1 (n_1557), .A2 (n_1414), .B1 (n_1412), .B2 (n_1410));
OAI21_X1 i_1204 (.ZN (n_4876), .A (n_1403), .B1 (n_1409), .B2 (n_1401));
OAI21_X1 i_1203 (.ZN (n_4867), .A (n_1397), .B1 (n_1399), .B2 (n_1395));
AOI21_X1 i_1202 (.ZN (n_1333), .A (n_4924), .B1 (n_4923), .B2 (n_1392));
INV_X1 i_1200 (.ZN (n_4927), .A (n_1333));
AOI21_X1 i_1199 (.ZN (n_4918), .A (n_1455), .B1 (n_1450), .B2 (n_1434));
AOI21_X1 i_1198 (.ZN (n_1332), .A (n_1361), .B1 (inputB[14]), .B2 (inputA[27]));
INV_X1 i_1196 (.ZN (n_1331), .A (n_1332));
NAND3_X1 i_1195 (.ZN (n_1329), .A1 (inputB[14]), .A2 (inputA[27]), .A3 (n_1361));
NAND2_X1 i_1194 (.ZN (n_1328), .A1 (n_1331), .A2 (n_1329));
NAND2_X1 i_1192 (.ZN (n_1324), .A1 (inputB[16]), .A2 (inputA[25]));
XOR2_X1 i_1191 (.Z (n_5031), .A (n_1328), .B (n_1324));
AND2_X1 i_1190 (.ZN (n_1319), .A1 (inputB[17]), .A2 (inputA[24]));
AOI21_X1 i_1189 (.ZN (n_1318), .A (n_1319), .B1 (inputB[18]), .B2 (inputA[23]));
INV_X1 i_1188 (.ZN (n_1314), .A (n_1318));
NAND3_X1 i_1187 (.ZN (n_1309), .A1 (inputB[18]), .A2 (inputA[23]), .A3 (n_1319));
NAND2_X1 i_1186 (.ZN (n_1305), .A1 (n_1314), .A2 (n_1309));
NAND2_X1 i_1185 (.ZN (n_1304), .A1 (inputB[19]), .A2 (inputA[22]));
XOR2_X1 i_1184 (.Z (n_5024), .A (n_1305), .B (n_1304));
AOI22_X1 i_1183 (.ZN (n_1300), .A1 (inputB[24]), .A2 (inputA[17]), .B1 (inputB[23]), .B2 (inputA[18]));
INV_X1 i_1182 (.ZN (n_1299), .A (n_1300));
NAND2_X1 i_1181 (.ZN (n_1298), .A1 (inputB[24]), .A2 (inputA[18]));
INV_X1 i_1180 (.ZN (n_1297), .A (n_1298));
NAND3_X1 i_1179 (.ZN (n_1295), .A1 (inputB[23]), .A2 (inputA[17]), .A3 (n_1297));
NAND2_X1 i_1178 (.ZN (n_1294), .A1 (n_1299), .A2 (n_1295));
NAND2_X1 i_1177 (.ZN (n_1293), .A1 (inputB[25]), .A2 (inputA[16]));
XOR2_X1 i_1176 (.Z (n_5010), .A (n_1294), .B (n_1293));
NAND2_X1 i_1175 (.ZN (n_1292), .A1 (inputB[26]), .A2 (inputA[15]));
INV_X1 i_1174 (.ZN (n_1291), .A (n_1292));
NAND2_X1 i_1173 (.ZN (n_1290), .A1 (n_1404), .A2 (n_1291));
OAI21_X1 i_1172 (.ZN (n_1289), .A (n_1290), .B1 (n_1404), .B2 (n_1291));
NAND2_X1 i_1171 (.ZN (n_1288), .A1 (inputB[28]), .A2 (inputA[13]));
XOR2_X1 i_1170 (.Z (n_5003), .A (n_1289), .B (n_1288));
AOI21_X1 i_1169 (.ZN (n_1287), .A (n_4934), .B1 (n_4933), .B2 (n_1354));
INV_X1 i_1168 (.ZN (n_4937), .A (n_1287));
AOI21_X1 i_1167 (.ZN (n_1286), .A (n_4929), .B1 (n_4928), .B2 (n_1393));
INV_X1 i_1166 (.ZN (n_1285), .A (n_1286));
XNOR2_X1 i_1165 (.ZN (n_5055), .A (n_5053), .B (n_1286));
OAI21_X1 i_1164 (.ZN (n_1284), .A (n_1360), .B1 (n_1363), .B2 (n_1357));
XOR2_X1 i_1162 (.Z (n_5045), .A (n_5043), .B (n_1284));
AOI21_X1 i_1161 (.ZN (n_1281), .A (n_4944), .B1 (n_4943), .B2 (n_1367));
INV_X1 i_1160 (.ZN (n_4947), .A (n_1281));
AOI21_X1 i_1158 (.ZN (n_1280), .A (n_4949), .B1 (n_4948), .B2 (n_1347));
INV_X1 i_1157 (.ZN (n_4952), .A (n_1280));
NAND2_X1 i_1156 (.ZN (n_1279), .A1 (inputB[12]), .A2 (inputA[30]));
NAND3_X1 i_1154 (.ZN (n_1278), .A1 (inputB[12]), .A2 (inputA[30]), .A3 (n_1430));
AOI22_X1 i_1153 (.ZN (n_1277), .A1 (inputB[12]), .A2 (inputA[29]), .B1 (inputB[11]), .B2 (inputA[30]));
INV_X1 i_1152 (.ZN (n_1274), .A (n_1277));
NAND2_X1 i_1150 (.ZN (n_1273), .A1 (n_1278), .A2 (n_1274));
NAND2_X1 i_1149 (.ZN (n_1269), .A1 (inputB[13]), .A2 (inputA[28]));
XOR2_X1 i_1148 (.Z (n_1265), .A (n_1273), .B (n_1269));
XOR2_X1 i_1147 (.Z (n_5060), .A (n_5058), .B (n_1265));
AND2_X1 i_1146 (.ZN (n_1264), .A1 (inputB[31]), .A2 (inputA[10]));
AOI22_X1 i_1145 (.ZN (n_1263), .A1 (inputB[30]), .A2 (inputA[11]), .B1 (inputB[29]), .B2 (inputA[12]));
NAND2_X1 i_1144 (.ZN (n_1259), .A1 (inputB[30]), .A2 (inputA[12]));
INV_X1 i_1143 (.ZN (n_1255), .A (n_1259));
NAND3_X1 i_1142 (.ZN (n_1254), .A1 (inputB[29]), .A2 (inputA[11]), .A3 (n_1255));
INV_X1 i_1141 (.ZN (n_1250), .A (n_1254));
NOR2_X1 i_1140 (.ZN (n_1249), .A1 (n_1263), .A2 (n_1250));
XNOR2_X1 i_1139 (.ZN (n_1248), .A (n_1264), .B (n_1249));
XOR2_X1 i_1138 (.Z (n_5070), .A (n_5068), .B (n_1248));
NAND2_X1 i_1137 (.ZN (n_1247), .A1 (inputB[21]), .A2 (inputA[21]));
INV_X1 i_1136 (.ZN (n_1246), .A (n_1247));
NAND2_X1 i_1135 (.ZN (n_1243), .A1 (n_1413), .A2 (n_1246));
AOI22_X1 i_1134 (.ZN (n_1242), .A1 (inputB[21]), .A2 (inputA[20]), .B1 (inputB[20]), .B2 (inputA[21]));
INV_X1 i_1133 (.ZN (n_1241), .A (n_1242));
NAND2_X1 i_1132 (.ZN (n_1240), .A1 (n_1243), .A2 (n_1241));
NAND2_X1 i_1131 (.ZN (n_1237), .A1 (inputB[22]), .A2 (inputA[19]));
XOR2_X1 i_1130 (.Z (n_1236), .A (n_1240), .B (n_1237));
XOR2_X1 i_1128 (.Z (n_5065), .A (n_5063), .B (n_1236));
AOI21_X1 i_1127 (.ZN (n_1235), .A (n_4939), .B1 (n_4938), .B2 (n_1356));
INV_X1 i_1126 (.ZN (n_1234), .A (n_1235));
XNOR2_X1 i_1124 (.ZN (n_5080), .A (n_5078), .B (n_1235));
AOI21_X1 i_1123 (.ZN (n_1233), .A (n_1377), .B1 (n_1381), .B2 (n_1371));
XOR2_X1 i_1122 (.Z (n_1231), .A (n_5048), .B (n_1233));
XOR2_X1 i_1120 (.Z (n_5075), .A (n_5073), .B (n_1231));
AOI21_X1 i_1119 (.ZN (n_1230), .A (n_4969), .B1 (n_4968), .B2 (n_1342));
INV_X1 i_1118 (.ZN (n_4972), .A (n_1230));
AOI21_X1 i_1117 (.ZN (n_1229), .A (n_4954), .B1 (n_4953), .B2 (n_1350));
INV_X1 i_1116 (.ZN (n_1228), .A (n_1229));
XNOR2_X1 i_1115 (.ZN (n_5085), .A (n_5083), .B (n_1229));
AOI21_X1 i_1114 (.ZN (n_1227), .A (n_4959), .B1 (n_4958), .B2 (n_1353));
INV_X1 i_1113 (.ZN (n_1226), .A (n_1227));
XNOR2_X1 i_1112 (.ZN (n_5090), .A (n_5088), .B (n_1227));
AOI21_X1 i_1111 (.ZN (n_1225), .A (n_4979), .B1 (n_4978), .B2 (n_1337));
INV_X1 i_1110 (.ZN (n_4982), .A (n_1225));
AOI21_X1 i_1109 (.ZN (n_1223), .A (n_4974), .B1 (n_4973), .B2 (n_1340));
INV_X1 i_1108 (.ZN (n_1222), .A (n_1223));
XNOR2_X1 i_1107 (.ZN (n_5100), .A (n_5098), .B (n_1223));
AOI21_X1 i_1106 (.ZN (n_1218), .A (n_4851), .B1 (n_4850), .B2 (n_1465));
INV_X1 i_1105 (.ZN (n_1213), .A (n_1218));
AOI21_X1 i_1104 (.ZN (n_1212), .A (n_4984), .B1 (n_4983), .B2 (n_1213));
INV_X1 i_1103 (.ZN (n_4987), .A (n_1212));
OAI21_X1 i_1102 (.ZN (n_5039), .A (n_1278), .B1 (n_1277), .B2 (n_1269));
OAI21_X1 i_1101 (.ZN (n_5032), .A (n_1329), .B1 (n_1332), .B2 (n_1324));
OAI21_X1 i_1100 (.ZN (n_5018), .A (n_1243), .B1 (n_1242), .B2 (n_1237));
OAI21_X1 i_1099 (.ZN (n_5011), .A (n_1295), .B1 (n_1300), .B2 (n_1293));
AOI21_X1 i_1097 (.ZN (n_4995), .A (n_1263), .B1 (n_1264), .B2 (n_1254));
AOI21_X1 i_1096 (.ZN (n_1209), .A (n_5049), .B1 (n_5048), .B2 (n_1233));
INV_X1 i_1095 (.ZN (n_5052), .A (n_1209));
OAI211_X1 i_1093 (.ZN (n_1208), .A (inputB[13]), .B (inputA[29]), .C1 (n_5758), .C2 (n_5753));
AOI211_X1 i_1092 (.ZN (n_1204), .A (n_5758), .B (n_5753), .C1 (inputB[13]), .C2 (inputA[29]));
INV_X1 i_1091 (.ZN (n_1203), .A (n_1204));
NAND2_X1 i_1090 (.ZN (n_1202), .A1 (n_1208), .A2 (n_1203));
XOR2_X1 i_1089 (.Z (n_5157), .A (n_1279), .B (n_1202));
AND2_X1 i_1088 (.ZN (n_1201), .A1 (inputB[14]), .A2 (inputA[28]));
AOI21_X1 i_1087 (.ZN (n_1200), .A (n_1201), .B1 (inputB[15]), .B2 (inputA[27]));
INV_X1 i_1086 (.ZN (n_1199), .A (n_1200));
NAND3_X1 i_1085 (.ZN (n_1198), .A1 (inputB[15]), .A2 (inputA[27]), .A3 (n_1201));
NAND2_X1 i_1084 (.ZN (n_1197), .A1 (n_1199), .A2 (n_1198));
NAND2_X1 i_1083 (.ZN (n_1196), .A1 (inputB[16]), .A2 (inputA[26]));
XOR2_X1 i_1082 (.Z (n_5151), .A (n_1197), .B (n_1196));
NAND2_X1 i_1081 (.ZN (n_1195), .A1 (inputB[20]), .A2 (inputA[22]));
INV_X1 i_1080 (.ZN (n_1194), .A (n_1195));
NAND2_X1 i_1079 (.ZN (n_1193), .A1 (n_1246), .A2 (n_1194));
NAND2_X1 i_1078 (.ZN (n_1191), .A1 (n_1247), .A2 (n_1195));
AND2_X1 i_1077 (.ZN (n_1190), .A1 (n_1193), .A2 (n_1191));
AND2_X1 i_1076 (.ZN (n_1189), .A1 (inputB[22]), .A2 (inputA[20]));
XOR2_X1 i_1075 (.Z (n_5137), .A (n_1190), .B (n_1189));
NAND2_X1 i_1074 (.ZN (n_1188), .A1 (inputB[23]), .A2 (inputA[19]));
INV_X1 i_1073 (.ZN (n_1187), .A (n_1188));
NAND2_X1 i_1072 (.ZN (n_1185), .A1 (n_1297), .A2 (n_1187));
OAI21_X1 i_1070 (.ZN (n_1184), .A (n_1185), .B1 (n_1297), .B2 (n_1187));
NAND2_X1 i_1069 (.ZN (n_1183), .A1 (inputB[25]), .A2 (inputA[17]));
XOR2_X1 i_1068 (.Z (n_5130), .A (n_1184), .B (n_1183));
NAND2_X1 i_1066 (.ZN (n_1182), .A1 (inputB[29]), .A2 (inputA[13]));
INV_X1 i_1065 (.ZN (n_1181), .A (n_1182));
NAND2_X1 i_1064 (.ZN (n_1180), .A1 (n_1255), .A2 (n_1181));
NAND2_X1 i_1063 (.ZN (n_1177), .A1 (n_1259), .A2 (n_1182));
AND2_X1 i_1062 (.ZN (n_1176), .A1 (n_1180), .A2 (n_1177));
NAND2_X1 i_1061 (.ZN (n_1172), .A1 (inputB[31]), .A2 (inputA[11]));
XOR2_X1 i_1060 (.Z (n_5114), .A (n_1176), .B (n_1172));
AOI21_X1 i_1059 (.ZN (n_1167), .A (n_5054), .B1 (n_5053), .B2 (n_1285));
INV_X1 i_1058 (.ZN (n_5057), .A (n_1167));
OAI21_X1 i_1057 (.ZN (n_1162), .A (n_1309), .B1 (n_1318), .B2 (n_1304));
XOR2_X1 i_1056 (.Z (n_5166), .A (n_5164), .B (n_1162));
AOI21_X1 i_1055 (.ZN (n_1158), .A (n_5069), .B1 (n_5068), .B2 (n_1248));
INV_X1 i_1054 (.ZN (n_5072), .A (n_1158));
AOI21_X1 i_1053 (.ZN (n_1157), .A (n_5059), .B1 (n_5058), .B2 (n_1265));
INV_X1 i_1051 (.ZN (n_5062), .A (n_1157));
AOI21_X1 i_1050 (.ZN (n_1156), .A (n_5044), .B1 (n_5043), .B2 (n_1284));
INV_X1 i_1049 (.ZN (n_1155), .A (n_1156));
XNOR2_X1 i_1048 (.ZN (n_5176), .A (n_5174), .B (n_1156));
AOI21_X1 i_1047 (.ZN (n_1153), .A (n_5074), .B1 (n_5073), .B2 (n_1231));
INV_X1 i_1046 (.ZN (n_5077), .A (n_1153));
NAND2_X1 i_1045 (.ZN (n_1152), .A1 (inputB[27]), .A2 (inputA[16]));
INV_X1 i_1044 (.ZN (n_1151), .A (n_1152));
NAND2_X1 i_1043 (.ZN (n_1150), .A1 (n_1291), .A2 (n_1151));
AOI22_X1 i_1042 (.ZN (n_1149), .A1 (inputB[27]), .A2 (inputA[15]), .B1 (inputB[26]), .B2 (inputA[16]));
INV_X1 i_1041 (.ZN (n_1148), .A (n_1149));
NAND2_X1 i_1040 (.ZN (n_1146), .A1 (n_1150), .A2 (n_1148));
NAND2_X1 i_1039 (.ZN (n_1145), .A1 (inputB[28]), .A2 (inputA[14]));
XOR2_X1 i_1038 (.Z (n_1144), .A (n_1146), .B (n_1145));
XOR2_X1 i_1037 (.Z (n_5186), .A (n_5184), .B (n_1144));
AOI22_X1 i_1036 (.ZN (n_1143), .A1 (n_1405), .A2 (n_1292), .B1 (n_1290), .B2 (n_1288));
XOR2_X1 i_1035 (.Z (n_1142), .A (n_5169), .B (n_1143));
XOR2_X1 i_1034 (.Z (n_5191), .A (n_5189), .B (n_1142));
AOI21_X1 i_1033 (.ZN (n_1140), .A (n_5084), .B1 (n_5083), .B2 (n_1228));
INV_X1 i_1032 (.ZN (n_5087), .A (n_1140));
AOI21_X1 i_1031 (.ZN (n_1139), .A (n_5089), .B1 (n_5088), .B2 (n_1226));
INV_X1 i_1030 (.ZN (n_5092), .A (n_1139));
AOI21_X1 i_1029 (.ZN (n_1138), .A (n_5079), .B1 (n_5078), .B2 (n_1234));
INV_X1 i_1028 (.ZN (n_1134), .A (n_1138));
XNOR2_X1 i_1027 (.ZN (n_5201), .A (n_5199), .B (n_1138));
NAND2_X1 i_1026 (.ZN (n_1129), .A1 (inputB[18]), .A2 (inputA[25]));
NAND3_X1 i_1025 (.ZN (n_1125), .A1 (inputB[18]), .A2 (inputA[25]), .A3 (n_1319));
AOI22_X1 i_1024 (.ZN (n_1124), .A1 (inputB[18]), .A2 (inputA[24]), .B1 (inputB[17]), .B2 (inputA[25]));
INV_X1 i_1023 (.ZN (n_1123), .A (n_1124));
NAND2_X1 i_1022 (.ZN (n_1122), .A1 (n_1125), .A2 (n_1123));
NAND2_X1 i_1021 (.ZN (n_1121), .A1 (inputB[19]), .A2 (inputA[23]));
XOR2_X1 i_1020 (.Z (n_1120), .A (n_1122), .B (n_1121));
XOR2_X1 i_1019 (.Z (n_1119), .A (n_5179), .B (n_1120));
XOR2_X1 i_1018 (.Z (n_5206), .A (n_5204), .B (n_1119));
AOI21_X1 i_1017 (.ZN (n_1118), .A (n_5064), .B1 (n_5063), .B2 (n_1236));
INV_X1 i_1016 (.ZN (n_1117), .A (n_1118));
XNOR2_X1 i_1015 (.ZN (n_1116), .A (n_5194), .B (n_1118));
XOR2_X1 i_1014 (.Z (n_5211), .A (n_5209), .B (n_1116));
AOI21_X1 i_1013 (.ZN (n_1115), .A (n_4964), .B1 (n_4963), .B2 (n_1346));
INV_X1 i_1012 (.ZN (n_1112), .A (n_1115));
AOI21_X1 i_1011 (.ZN (n_1111), .A (n_5094), .B1 (n_5093), .B2 (n_1112));
INV_X1 i_1010 (.ZN (n_1110), .A (n_1111));
XNOR2_X1 i_1009 (.ZN (n_5216), .A (n_5214), .B (n_1111));
XNOR2_X1 i_1008 (.ZN (n_1109), .A (n_5093), .B (n_1115));
AOI21_X1 i_1007 (.ZN (n_1108), .A (n_5104), .B1 (n_5103), .B2 (n_1109));
INV_X1 i_1006 (.ZN (n_5107), .A (n_1108));
OAI21_X1 i_1005 (.ZN (n_5152), .A (n_1198), .B1 (n_1200), .B2 (n_1196));
OAI21_X1 i_1004 (.ZN (n_5145), .A (n_1125), .B1 (n_1124), .B2 (n_1121));
AOI22_X1 i_1003 (.ZN (n_5131), .A1 (n_1298), .A2 (n_1188), .B1 (n_1185), .B2 (n_1183));
OAI21_X1 i_1002 (.ZN (n_5124), .A (n_1150), .B1 (n_1149), .B2 (n_1145));
AOI21_X1 i_1001 (.ZN (n_1105), .A (n_5170), .B1 (n_5169), .B2 (n_1143));
INV_X1 i_1000 (.ZN (n_5173), .A (n_1105));
AOI21_X1 i_999 (.ZN (n_1104), .A (n_5165), .B1 (n_5164), .B2 (n_1162));
INV_X1 i_998 (.ZN (n_5168), .A (n_1104));
NAND2_X1 i_997 (.ZN (n_1100), .A1 (inputB[15]), .A2 (inputA[29]));
INV_X1 i_996 (.ZN (n_1096), .A (n_1100));
NAND2_X1 i_995 (.ZN (n_1095), .A1 (n_1201), .A2 (n_1096));
AOI22_X1 i_994 (.ZN (n_1094), .A1 (inputB[15]), .A2 (inputA[28]), .B1 (inputB[14]), .B2 (inputA[29]));
INV_X1 i_993 (.ZN (n_1093), .A (n_1094));
NAND2_X1 i_992 (.ZN (n_1091), .A1 (n_1095), .A2 (n_1093));
NAND2_X1 i_991 (.ZN (n_1090), .A1 (inputB[16]), .A2 (inputA[27]));
XOR2_X1 i_990 (.Z (n_5267), .A (n_1091), .B (n_1090));
NAND2_X1 i_989 (.ZN (n_1089), .A1 (inputB[17]), .A2 (inputA[26]));
OR2_X1 i_988 (.ZN (n_1088), .A1 (n_1129), .A2 (n_1089));
NAND2_X1 i_987 (.ZN (n_1087), .A1 (n_1129), .A2 (n_1089));
AND2_X1 i_986 (.ZN (n_1086), .A1 (n_1088), .A2 (n_1087));
AND2_X1 i_985 (.ZN (n_1085), .A1 (inputB[19]), .A2 (inputA[24]));
XOR2_X1 i_984 (.Z (n_5260), .A (n_1086), .B (n_1085));
AOI22_X1 i_983 (.ZN (n_1083), .A1 (inputB[24]), .A2 (inputA[19]), .B1 (inputB[23]), .B2 (inputA[20]));
INV_X1 i_982 (.ZN (n_1082), .A (n_1083));
NAND2_X1 i_981 (.ZN (n_1081), .A1 (inputB[24]), .A2 (inputA[20]));
INV_X1 i_980 (.ZN (n_1080), .A (n_1081));
NAND2_X1 i_979 (.ZN (n_1079), .A1 (n_1187), .A2 (n_1080));
NAND2_X1 i_978 (.ZN (n_1076), .A1 (n_1082), .A2 (n_1079));
NAND2_X1 i_977 (.ZN (n_1075), .A1 (inputB[25]), .A2 (inputA[18]));
XOR2_X1 i_976 (.Z (n_5246), .A (n_1076), .B (n_1075));
NAND2_X1 i_975 (.ZN (n_1071), .A1 (inputB[26]), .A2 (inputA[17]));
INV_X1 i_974 (.ZN (n_1067), .A (n_1071));
NAND2_X1 i_973 (.ZN (n_1066), .A1 (n_1151), .A2 (n_1067));
NAND2_X1 i_972 (.ZN (n_1065), .A1 (n_1152), .A2 (n_1071));
AND2_X1 i_971 (.ZN (n_1064), .A1 (n_1066), .A2 (n_1065));
AND2_X1 i_970 (.ZN (n_1063), .A1 (inputB[28]), .A2 (inputA[15]));
XOR2_X1 i_969 (.Z (n_5239), .A (n_1064), .B (n_1063));
AOI21_X1 i_968 (.ZN (n_1062), .A (n_5175), .B1 (n_5174), .B2 (n_1155));
INV_X1 i_967 (.ZN (n_5178), .A (n_1062));
NAND2_X1 i_966 (.ZN (n_1061), .A1 (n_1177), .A2 (n_1172));
NAND2_X1 i_965 (.ZN (n_1060), .A1 (n_1180), .A2 (n_1061));
XOR2_X1 i_964 (.Z (n_5287), .A (n_5285), .B (n_1060));
AOI21_X1 i_963 (.ZN (n_1059), .A (n_5185), .B1 (n_5184), .B2 (n_1144));
INV_X1 i_962 (.ZN (n_5188), .A (n_1059));
AOI21_X1 i_961 (.ZN (n_1058), .A (n_5180), .B1 (n_5179), .B2 (n_1120));
INV_X1 i_960 (.ZN (n_5183), .A (n_1058));
AOI21_X1 i_959 (.ZN (n_1057), .A (n_5195), .B1 (n_5194), .B2 (n_1117));
INV_X1 i_958 (.ZN (n_5198), .A (n_1057));
AOI21_X1 i_957 (.ZN (n_1055), .A (n_5190), .B1 (n_5189), .B2 (n_1142));
INV_X1 i_956 (.ZN (n_5193), .A (n_1055));
AND2_X1 i_955 (.ZN (n_1054), .A1 (inputB[21]), .A2 (inputA[23]));
NAND2_X1 i_954 (.ZN (n_1051), .A1 (n_1194), .A2 (n_1054));
AOI22_X1 i_953 (.ZN (n_1050), .A1 (inputB[21]), .A2 (inputA[22]), .B1 (inputB[20]), .B2 (inputA[23]));
INV_X1 i_952 (.ZN (n_1049), .A (n_1050));
NAND2_X1 i_951 (.ZN (n_1048), .A1 (n_1051), .A2 (n_1049));
NAND2_X1 i_950 (.ZN (n_1047), .A1 (inputB[22]), .A2 (inputA[21]));
XOR2_X1 i_949 (.Z (n_1044), .A (n_1048), .B (n_1047));
XOR2_X1 i_948 (.Z (n_5297), .A (n_5295), .B (n_1044));
AOI21_X1 i_947 (.ZN (n_1043), .A (n_5200), .B1 (n_5199), .B2 (n_1134));
INV_X1 i_946 (.ZN (n_5203), .A (n_1043));
NAND2_X1 i_945 (.ZN (n_1042), .A1 (n_1191), .A2 (n_1189));
NAND2_X1 i_944 (.ZN (n_1041), .A1 (n_1193), .A2 (n_1042));
XOR2_X1 i_943 (.Z (n_1038), .A (n_5280), .B (n_1041));
XOR2_X1 i_942 (.Z (n_5307), .A (n_5305), .B (n_1038));
AOI21_X1 i_941 (.ZN (n_1037), .A (n_5205), .B1 (n_5204), .B2 (n_1119));
INV_X1 i_940 (.ZN (n_5208), .A (n_1037));
AOI21_X1 i_939 (.ZN (n_1036), .A (n_5210), .B1 (n_5209), .B2 (n_1116));
INV_X1 i_938 (.ZN (n_5213), .A (n_1036));
NAND2_X1 i_937 (.ZN (n_1035), .A1 (inputB[12]), .A2 (inputA[31]));
AND2_X1 i_936 (.ZN (n_1033), .A1 (inputB[13]), .A2 (inputA[30]));
NAND2_X1 i_935 (.ZN (n_1032), .A1 (n_1035), .A2 (n_1033));
OAI21_X1 i_934 (.ZN (n_1031), .A (n_1032), .B1 (n_1035), .B2 (n_1033));
AOI21_X1 i_933 (.ZN (n_1028), .A (n_1204), .B1 (n_1279), .B2 (n_1208));
INV_X1 i_932 (.ZN (n_1027), .A (n_1028));
XNOR2_X1 i_931 (.ZN (n_1026), .A (n_1031), .B (n_1028));
XOR2_X1 i_930 (.Z (n_1025), .A (n_5290), .B (n_1026));
XOR2_X1 i_929 (.Z (n_1024), .A (n_5310), .B (n_1025));
XOR2_X1 i_928 (.Z (n_5322), .A (n_5320), .B (n_1024));
NAND2_X1 i_927 (.ZN (n_1023), .A1 (inputB[30]), .A2 (inputA[14]));
INV_X1 i_926 (.ZN (n_1021), .A (n_1023));
AOI22_X1 i_925 (.ZN (n_1020), .A1 (inputB[30]), .A2 (inputA[13]), .B1 (inputB[29]), .B2 (inputA[14]));
AOI21_X1 i_924 (.ZN (n_1019), .A (n_1020), .B1 (n_1181), .B2 (n_1021));
NAND2_X1 i_923 (.ZN (n_1018), .A1 (inputB[31]), .A2 (inputA[12]));
XOR2_X1 i_922 (.Z (n_1017), .A (n_1019), .B (n_1018));
XOR2_X1 i_921 (.Z (n_1016), .A (n_5300), .B (n_1017));
XOR2_X1 i_920 (.Z (n_1015), .A (n_5315), .B (n_1016));
XOR2_X1 i_919 (.Z (n_5327), .A (n_5325), .B (n_1015));
AOI21_X1 i_918 (.ZN (n_1014), .A (n_5099), .B1 (n_5098), .B2 (n_1222));
INV_X1 i_917 (.ZN (n_1013), .A (n_1014));
AOI21_X1 i_916 (.ZN (n_1012), .A (n_5220), .B1 (n_5219), .B2 (n_1013));
INV_X1 i_915 (.ZN (n_5223), .A (n_1012));
NAND2_X1 i_914 (.ZN (n_447), .A1 (inputB[13]), .A2 (inputA[31]));
OAI21_X1 i_913 (.ZN (n_5268), .A (n_1095), .B1 (n_1094), .B2 (n_1090));
OAI21_X1 i_912 (.ZN (n_5254), .A (n_1051), .B1 (n_1050), .B2 (n_1047));
OAI21_X1 i_911 (.ZN (n_5247), .A (n_1079), .B1 (n_1083), .B2 (n_1075));
AOI22_X1 i_910 (.ZN (n_1011), .A1 (n_1181), .A2 (n_1021), .B1 (n_1019), .B2 (n_1018));
INV_X1 i_909 (.ZN (n_5231), .A (n_1011));
AOI21_X1 i_908 (.ZN (n_1010), .A (n_5286), .B1 (n_5285), .B2 (n_1060));
INV_X1 i_907 (.ZN (n_5289), .A (n_1010));
OAI21_X1 i_906 (.ZN (n_5275), .A (n_1032), .B1 (n_1031), .B2 (n_1027));
NAND3_X1 i_905 (.ZN (n_1009), .A1 (inputB[14]), .A2 (inputA[30]), .A3 (n_1096));
INV_X1 i_904 (.ZN (n_1008), .A (n_1009));
AOI21_X1 i_903 (.ZN (n_1007), .A (n_1096), .B1 (inputB[14]), .B2 (inputA[30]));
NOR2_X1 i_902 (.ZN (n_1006), .A1 (n_1008), .A2 (n_1007));
NAND2_X1 i_901 (.ZN (n_1005), .A1 (inputB[16]), .A2 (inputA[28]));
XNOR2_X1 i_900 (.ZN (n_5378), .A (n_1006), .B (n_1005));
AOI21_X1 i_899 (.ZN (n_1004), .A (n_1054), .B1 (inputB[20]), .B2 (inputA[24]));
INV_X1 i_898 (.ZN (n_1003), .A (n_1004));
NAND3_X1 i_897 (.ZN (n_1002), .A1 (inputB[20]), .A2 (inputA[24]), .A3 (n_1054));
NAND2_X1 i_896 (.ZN (n_1001), .A1 (n_1003), .A2 (n_1002));
NAND2_X1 i_895 (.ZN (n_1000), .A1 (inputB[22]), .A2 (inputA[22]));
XOR2_X1 i_894 (.Z (n_5364), .A (n_1001), .B (n_1000));
NAND2_X1 i_893 (.ZN (n_999), .A1 (inputB[23]), .A2 (inputA[21]));
INV_X1 i_892 (.ZN (n_998), .A (n_999));
NAND2_X1 i_891 (.ZN (n_997), .A1 (n_1080), .A2 (n_998));
OAI21_X1 i_890 (.ZN (n_996), .A (n_997), .B1 (n_1080), .B2 (n_998));
NAND2_X1 i_889 (.ZN (n_995), .A1 (inputB[25]), .A2 (inputA[19]));
XOR2_X1 i_888 (.Z (n_5357), .A (n_996), .B (n_995));
NAND2_X1 i_887 (.ZN (n_994), .A1 (inputB[29]), .A2 (inputA[15]));
INV_X1 i_886 (.ZN (n_993), .A (n_994));
NAND2_X1 i_885 (.ZN (n_992), .A1 (n_1021), .A2 (n_993));
NAND2_X1 i_884 (.ZN (n_990), .A1 (n_1023), .A2 (n_994));
AND2_X1 i_883 (.ZN (n_989), .A1 (n_992), .A2 (n_990));
NAND2_X1 i_882 (.ZN (n_988), .A1 (inputB[31]), .A2 (inputA[13]));
XOR2_X1 i_881 (.Z (n_5341), .A (n_989), .B (n_988));
NAND2_X1 i_880 (.ZN (n_987), .A1 (n_1065), .A2 (n_1063));
NAND2_X1 i_879 (.ZN (n_986), .A1 (n_1066), .A2 (n_987));
XOR2_X1 i_878 (.Z (n_5390), .A (n_5388), .B (n_986));
AOI21_X1 i_877 (.ZN (n_985), .A (n_5301), .B1 (n_5300), .B2 (n_1017));
INV_X1 i_876 (.ZN (n_5304), .A (n_985));
AOI21_X1 i_875 (.ZN (n_984), .A (n_5296), .B1 (n_5295), .B2 (n_1044));
INV_X1 i_874 (.ZN (n_5299), .A (n_984));
AOI21_X1 i_873 (.ZN (n_983), .A (n_5281), .B1 (n_5280), .B2 (n_1041));
INV_X1 i_872 (.ZN (n_982), .A (n_983));
XNOR2_X1 i_871 (.ZN (n_5395), .A (n_5393), .B (n_983));
AOI21_X1 i_870 (.ZN (n_981), .A (n_5306), .B1 (n_5305), .B2 (n_1038));
INV_X1 i_869 (.ZN (n_5309), .A (n_981));
NAND2_X1 i_868 (.ZN (n_980), .A1 (inputB[18]), .A2 (inputA[27]));
OR2_X1 i_867 (.ZN (n_979), .A1 (n_1089), .A2 (n_980));
AOI22_X1 i_866 (.ZN (n_978), .A1 (inputB[18]), .A2 (inputA[26]), .B1 (inputB[17]), .B2 (inputA[27]));
INV_X1 i_865 (.ZN (n_977), .A (n_978));
NAND2_X1 i_864 (.ZN (n_976), .A1 (n_979), .A2 (n_977));
NAND2_X1 i_863 (.ZN (n_975), .A1 (inputB[19]), .A2 (inputA[25]));
XOR2_X1 i_862 (.Z (n_974), .A (n_976), .B (n_975));
XOR2_X1 i_861 (.Z (n_5400), .A (n_5398), .B (n_974));
AOI21_X1 i_860 (.ZN (n_973), .A (n_5311), .B1 (n_5310), .B2 (n_1025));
INV_X1 i_859 (.ZN (n_5314), .A (n_973));
NAND2_X1 i_858 (.ZN (n_972), .A1 (n_1087), .A2 (n_1085));
NAND2_X1 i_857 (.ZN (n_971), .A1 (n_1088), .A2 (n_972));
XOR2_X1 i_856 (.Z (n_970), .A (n_5383), .B (n_971));
XOR2_X1 i_855 (.Z (n_5410), .A (n_5408), .B (n_970));
AOI21_X1 i_854 (.ZN (n_969), .A (n_5316), .B1 (n_5315), .B2 (n_1016));
INV_X1 i_853 (.ZN (n_5319), .A (n_969));
AOI21_X1 i_852 (.ZN (n_968), .A (n_5321), .B1 (n_5320), .B2 (n_1024));
INV_X1 i_851 (.ZN (n_5324), .A (n_968));
AOI21_X1 i_850 (.ZN (n_967), .A (n_5291), .B1 (n_5290), .B2 (n_1026));
INV_X1 i_849 (.ZN (n_966), .A (n_967));
XNOR2_X1 i_848 (.ZN (n_965), .A (n_5413), .B (n_967));
XOR2_X1 i_847 (.Z (n_5425), .A (n_5423), .B (n_965));
NAND2_X1 i_846 (.ZN (n_964), .A1 (inputB[27]), .A2 (inputA[18]));
INV_X1 i_845 (.ZN (n_963), .A (n_964));
NAND2_X1 i_844 (.ZN (n_962), .A1 (n_1067), .A2 (n_963));
AOI22_X1 i_843 (.ZN (n_961), .A1 (inputB[27]), .A2 (inputA[17]), .B1 (inputB[26]), .B2 (inputA[18]));
INV_X1 i_842 (.ZN (n_960), .A (n_961));
NAND2_X1 i_841 (.ZN (n_959), .A1 (n_962), .A2 (n_960));
NAND2_X1 i_840 (.ZN (n_958), .A1 (inputB[28]), .A2 (inputA[16]));
XOR2_X1 i_839 (.Z (n_957), .A (n_959), .B (n_958));
XOR2_X1 i_838 (.Z (n_956), .A (n_5403), .B (n_957));
XOR2_X1 i_837 (.Z (n_955), .A (n_5418), .B (n_956));
XOR2_X1 i_836 (.Z (n_5430), .A (n_5428), .B (n_955));
AOI21_X1 i_835 (.ZN (n_954), .A (n_5215), .B1 (n_5214), .B2 (n_1110));
INV_X1 i_834 (.ZN (n_953), .A (n_954));
AOI21_X1 i_833 (.ZN (n_952), .A (n_5331), .B1 (n_5330), .B2 (n_953));
INV_X1 i_832 (.ZN (n_5334), .A (n_952));
OAI21_X1 i_831 (.ZN (n_5379), .A (n_1009), .B1 (n_1007), .B2 (n_1005));
OAI21_X1 i_830 (.ZN (n_5372), .A (n_979), .B1 (n_978), .B2 (n_975));
AOI22_X1 i_829 (.ZN (n_5358), .A1 (n_1081), .A2 (n_999), .B1 (n_997), .B2 (n_995));
OAI21_X1 i_828 (.ZN (n_5351), .A (n_962), .B1 (n_961), .B2 (n_958));
AOI21_X1 i_827 (.ZN (n_951), .A (n_5389), .B1 (n_5388), .B2 (n_986));
INV_X1 i_826 (.ZN (n_5392), .A (n_951));
AOI21_X1 i_825 (.ZN (n_950), .A (n_5384), .B1 (n_5383), .B2 (n_971));
INV_X1 i_824 (.ZN (n_5387), .A (n_950));
NAND2_X1 i_823 (.ZN (n_949), .A1 (inputB[17]), .A2 (inputA[28]));
OR2_X1 i_822 (.ZN (n_948), .A1 (n_980), .A2 (n_949));
NAND2_X1 i_821 (.ZN (n_947), .A1 (n_980), .A2 (n_949));
AND2_X1 i_820 (.ZN (n_946), .A1 (n_948), .A2 (n_947));
AND2_X1 i_819 (.ZN (n_945), .A1 (inputB[19]), .A2 (inputA[26]));
XOR2_X1 i_818 (.Z (n_5474), .A (n_946), .B (n_945));
AND2_X1 i_817 (.ZN (n_944), .A1 (inputB[20]), .A2 (inputA[25]));
AOI21_X1 i_816 (.ZN (n_943), .A (n_944), .B1 (inputB[21]), .B2 (inputA[24]));
INV_X1 i_815 (.ZN (n_942), .A (n_943));
NAND3_X1 i_814 (.ZN (n_941), .A1 (inputB[21]), .A2 (inputA[24]), .A3 (n_944));
NAND2_X1 i_813 (.ZN (n_940), .A1 (n_942), .A2 (n_941));
NAND2_X1 i_812 (.ZN (n_939), .A1 (inputB[22]), .A2 (inputA[23]));
XOR2_X1 i_811 (.Z (n_5467), .A (n_940), .B (n_939));
NAND2_X1 i_810 (.ZN (n_938), .A1 (inputB[26]), .A2 (inputA[19]));
INV_X1 i_809 (.ZN (n_937), .A (n_938));
NAND2_X1 i_808 (.ZN (n_936), .A1 (n_963), .A2 (n_937));
NAND2_X1 i_807 (.ZN (n_935), .A1 (n_964), .A2 (n_938));
AND2_X1 i_806 (.ZN (n_934), .A1 (n_936), .A2 (n_935));
AND2_X1 i_805 (.ZN (n_933), .A1 (inputB[28]), .A2 (inputA[17]));
XOR2_X1 i_804 (.Z (n_5453), .A (n_934), .B (n_933));
NAND2_X1 i_803 (.ZN (n_932), .A1 (inputB[30]), .A2 (inputA[16]));
INV_X1 i_802 (.ZN (n_931), .A (n_932));
AOI22_X1 i_801 (.ZN (n_930), .A1 (inputB[30]), .A2 (inputA[15]), .B1 (inputB[29]), .B2 (inputA[16]));
AOI21_X1 i_800 (.ZN (n_929), .A (n_930), .B1 (n_993), .B2 (n_931));
NAND2_X1 i_799 (.ZN (n_928), .A1 (inputB[31]), .A2 (inputA[14]));
XOR2_X1 i_798 (.Z (n_5444), .A (n_929), .B (n_928));
NAND2_X1 i_797 (.ZN (n_926), .A1 (n_990), .A2 (n_988));
NAND2_X1 i_796 (.ZN (n_925), .A1 (n_992), .A2 (n_926));
XOR2_X1 i_795 (.Z (n_5494), .A (n_5492), .B (n_925));
OAI21_X1 i_794 (.ZN (n_924), .A (n_1002), .B1 (n_1004), .B2 (n_1000));
XOR2_X1 i_793 (.Z (n_5489), .A (n_5487), .B (n_924));
AOI21_X1 i_792 (.ZN (n_923), .A (n_5399), .B1 (n_5398), .B2 (n_974));
INV_X1 i_791 (.ZN (n_5402), .A (n_923));
NAND2_X1 i_790 (.ZN (n_922), .A1 (inputB[16]), .A2 (inputA[30]));
NOR2_X1 i_789 (.ZN (n_921), .A1 (n_1100), .A2 (n_922));
AOI22_X1 i_788 (.ZN (n_920), .A1 (inputB[15]), .A2 (inputA[30]), .B1 (inputB[16]), .B2 (inputA[29]));
INV_X1 i_787 (.ZN (n_919), .A (n_920));
NOR2_X1 i_786 (.ZN (n_918), .A1 (n_921), .A2 (n_920));
NAND2_X1 i_785 (.ZN (n_917), .A1 (inputB[14]), .A2 (inputA[31]));
XOR2_X1 i_784 (.Z (n_916), .A (n_918), .B (n_917));
XOR2_X1 i_783 (.Z (n_5499), .A (n_5497), .B (n_916));
AOI21_X1 i_782 (.ZN (n_915), .A (n_5409), .B1 (n_5408), .B2 (n_970));
INV_X1 i_781 (.ZN (n_5412), .A (n_915));
AOI21_X1 i_780 (.ZN (n_914), .A (n_5394), .B1 (n_5393), .B2 (n_982));
INV_X1 i_779 (.ZN (n_913), .A (n_914));
XNOR2_X1 i_778 (.ZN (n_5509), .A (n_5507), .B (n_914));
AOI21_X1 i_777 (.ZN (n_912), .A (n_5404), .B1 (n_5403), .B2 (n_957));
INV_X1 i_776 (.ZN (n_911), .A (n_912));
XNOR2_X1 i_775 (.ZN (n_5514), .A (n_5512), .B (n_912));
AOI21_X1 i_774 (.ZN (n_910), .A (n_5419), .B1 (n_5418), .B2 (n_956));
INV_X1 i_773 (.ZN (n_5422), .A (n_910));
AOI21_X1 i_772 (.ZN (n_909), .A (n_5424), .B1 (n_5423), .B2 (n_965));
INV_X1 i_771 (.ZN (n_5427), .A (n_909));
AND2_X1 i_770 (.ZN (n_908), .A1 (inputB[24]), .A2 (inputA[22]));
NAND2_X1 i_769 (.ZN (n_907), .A1 (n_998), .A2 (n_908));
AOI22_X1 i_768 (.ZN (n_906), .A1 (inputB[24]), .A2 (inputA[21]), .B1 (inputB[23]), .B2 (inputA[22]));
INV_X1 i_767 (.ZN (n_905), .A (n_906));
NAND2_X1 i_766 (.ZN (n_904), .A1 (n_907), .A2 (n_905));
NAND2_X1 i_765 (.ZN (n_903), .A1 (inputB[25]), .A2 (inputA[20]));
XOR2_X1 i_764 (.Z (n_902), .A (n_904), .B (n_903));
XOR2_X1 i_763 (.Z (n_901), .A (n_5502), .B (n_902));
XOR2_X1 i_762 (.Z (n_5524), .A (n_5522), .B (n_901));
AOI21_X1 i_761 (.ZN (n_900), .A (n_5414), .B1 (n_5413), .B2 (n_966));
INV_X1 i_760 (.ZN (n_899), .A (n_900));
XNOR2_X1 i_759 (.ZN (n_898), .A (n_5517), .B (n_900));
XOR2_X1 i_758 (.Z (n_5529), .A (n_5527), .B (n_898));
AOI21_X1 i_757 (.ZN (n_897), .A (n_5326), .B1 (n_5325), .B2 (n_1015));
INV_X1 i_756 (.ZN (n_896), .A (n_897));
AOI21_X1 i_755 (.ZN (n_895), .A (n_5434), .B1 (n_5433), .B2 (n_896));
INV_X1 i_754 (.ZN (n_5437), .A (n_895));
NAND2_X1 i_753 (.ZN (n_894), .A1 (n_947), .A2 (n_945));
NAND2_X1 i_752 (.ZN (n_5475), .A1 (n_948), .A2 (n_894));
OAI21_X1 i_751 (.ZN (n_5468), .A (n_941), .B1 (n_943), .B2 (n_939));
NAND2_X1 i_750 (.ZN (n_893), .A1 (n_935), .A2 (n_933));
NAND2_X1 i_749 (.ZN (n_5454), .A1 (n_936), .A2 (n_893));
AOI22_X1 i_748 (.ZN (n_892), .A1 (n_993), .A2 (n_931), .B1 (n_929), .B2 (n_928));
INV_X1 i_747 (.ZN (n_5445), .A (n_892));
AOI21_X1 i_746 (.ZN (n_891), .A (n_5488), .B1 (n_5487), .B2 (n_924));
INV_X1 i_745 (.ZN (n_5491), .A (n_891));
AOI21_X1 i_744 (.ZN (n_890), .A (n_922), .B1 (inputB[15]), .B2 (inputA[31]));
INV_X1 i_743 (.ZN (n_889), .A (n_890));
AND3_X1 i_742 (.ZN (n_888), .A1 (inputB[15]), .A2 (inputA[31]), .A3 (n_922));
NOR2_X1 i_741 (.ZN (n_887), .A1 (n_890), .A2 (n_888));
AOI21_X1 i_740 (.ZN (n_886), .A (n_921), .B1 (n_919), .B2 (n_917));
XNOR2_X1 i_739 (.ZN (n_5580), .A (n_887), .B (n_886));
AOI22_X1 i_738 (.ZN (n_885), .A1 (inputB[21]), .A2 (inputA[25]), .B1 (inputB[20]), .B2 (inputA[26]));
INV_X1 i_737 (.ZN (n_884), .A (n_885));
NAND2_X1 i_736 (.ZN (n_883), .A1 (inputB[21]), .A2 (inputA[26]));
INV_X1 i_735 (.ZN (n_882), .A (n_883));
NAND2_X1 i_734 (.ZN (n_881), .A1 (n_944), .A2 (n_882));
NAND2_X1 i_733 (.ZN (n_880), .A1 (n_884), .A2 (n_881));
NAND2_X1 i_732 (.ZN (n_879), .A1 (inputB[22]), .A2 (inputA[24]));
XOR2_X1 i_731 (.Z (n_5566), .A (n_880), .B (n_879));
AOI21_X1 i_730 (.ZN (n_878), .A (n_908), .B1 (inputB[23]), .B2 (inputA[23]));
INV_X1 i_729 (.ZN (n_877), .A (n_878));
NAND3_X1 i_728 (.ZN (n_876), .A1 (inputB[23]), .A2 (inputA[23]), .A3 (n_908));
NAND2_X1 i_727 (.ZN (n_875), .A1 (n_877), .A2 (n_876));
NAND2_X1 i_726 (.ZN (n_874), .A1 (inputB[25]), .A2 (inputA[21]));
XOR2_X1 i_725 (.Z (n_5559), .A (n_875), .B (n_874));
NAND2_X1 i_724 (.ZN (n_873), .A1 (inputB[29]), .A2 (inputA[17]));
INV_X1 i_723 (.ZN (n_872), .A (n_873));
NAND2_X1 i_722 (.ZN (n_871), .A1 (n_931), .A2 (n_872));
NAND2_X1 i_721 (.ZN (n_870), .A1 (n_932), .A2 (n_873));
NAND2_X1 i_720 (.ZN (n_869), .A1 (n_871), .A2 (n_870));
NAND2_X1 i_719 (.ZN (n_868), .A1 (inputB[31]), .A2 (inputA[15]));
NAND2_X1 i_718 (.ZN (n_867), .A1 (n_870), .A2 (n_868));
XNOR2_X1 i_717 (.ZN (n_5543), .A (n_869), .B (n_868));
AOI21_X1 i_716 (.ZN (n_866), .A (n_5493), .B1 (n_5492), .B2 (n_925));
INV_X1 i_715 (.ZN (n_865), .A (n_866));
XNOR2_X1 i_714 (.ZN (n_5593), .A (n_5591), .B (n_866));
AOI21_X1 i_713 (.ZN (n_864), .A (n_5503), .B1 (n_5502), .B2 (n_902));
INV_X1 i_712 (.ZN (n_5506), .A (n_864));
AOI21_X1 i_711 (.ZN (n_863), .A (n_5498), .B1 (n_5497), .B2 (n_916));
INV_X1 i_710 (.ZN (n_5501), .A (n_863));
AOI21_X1 i_709 (.ZN (n_862), .A (n_5513), .B1 (n_5512), .B2 (n_911));
INV_X1 i_708 (.ZN (n_5516), .A (n_862));
AOI22_X1 i_707 (.ZN (n_861), .A1 (inputB[27]), .A2 (inputA[19]), .B1 (inputB[26]), .B2 (inputA[20]));
INV_X1 i_706 (.ZN (n_860), .A (n_861));
NAND3_X1 i_705 (.ZN (n_859), .A1 (inputB[27]), .A2 (inputA[20]), .A3 (n_937));
NAND2_X1 i_704 (.ZN (n_858), .A1 (n_860), .A2 (n_859));
NAND2_X1 i_703 (.ZN (n_857), .A1 (inputB[28]), .A2 (inputA[18]));
XOR2_X1 i_702 (.Z (n_856), .A (n_858), .B (n_857));
XOR2_X1 i_701 (.Z (n_5603), .A (n_5601), .B (n_856));
AOI21_X1 i_700 (.ZN (n_855), .A (n_5518), .B1 (n_5517), .B2 (n_899));
INV_X1 i_699 (.ZN (n_5521), .A (n_855));
AOI21_X1 i_698 (.ZN (n_854), .A (n_5508), .B1 (n_5507), .B2 (n_913));
INV_X1 i_697 (.ZN (n_853), .A (n_854));
XNOR2_X1 i_696 (.ZN (n_5613), .A (n_5611), .B (n_854));
AOI21_X1 i_695 (.ZN (n_852), .A (n_5523), .B1 (n_5522), .B2 (n_901));
INV_X1 i_694 (.ZN (n_5526), .A (n_852));
NAND2_X1 i_693 (.ZN (n_851), .A1 (inputB[18]), .A2 (inputA[29]));
OR2_X1 i_692 (.ZN (n_850), .A1 (n_949), .A2 (n_851));
AOI22_X1 i_691 (.ZN (n_849), .A1 (inputB[18]), .A2 (inputA[28]), .B1 (inputB[17]), .B2 (inputA[29]));
INV_X1 i_690 (.ZN (n_848), .A (n_849));
NAND2_X1 i_689 (.ZN (n_847), .A1 (n_850), .A2 (n_848));
NAND2_X1 i_688 (.ZN (n_846), .A1 (inputB[19]), .A2 (inputA[27]));
XOR2_X1 i_687 (.Z (n_845), .A (n_847), .B (n_846));
XOR2_X1 i_686 (.Z (n_844), .A (n_5596), .B (n_845));
XOR2_X1 i_685 (.Z (n_5618), .A (n_5616), .B (n_844));
AOI21_X1 i_684 (.ZN (n_843), .A (n_906), .B1 (n_907), .B2 (n_903));
XOR2_X1 i_683 (.Z (n_842), .A (n_5586), .B (n_843));
XOR2_X1 i_682 (.Z (n_841), .A (n_5606), .B (n_842));
XOR2_X1 i_681 (.Z (n_5623), .A (n_5621), .B (n_841));
AOI21_X1 i_680 (.ZN (n_840), .A (n_5429), .B1 (n_5428), .B2 (n_955));
INV_X1 i_679 (.ZN (n_839), .A (n_840));
AOI21_X1 i_678 (.ZN (n_838), .A (n_5533), .B1 (n_5532), .B2 (n_839));
INV_X1 i_677 (.ZN (n_5536), .A (n_838));
NAND2_X1 i_676 (.ZN (n_543), .A1 (inputB[16]), .A2 (inputA[31]));
OAI21_X1 i_675 (.ZN (n_5574), .A (n_850), .B1 (n_849), .B2 (n_846));
OAI21_X1 i_674 (.ZN (n_5560), .A (n_876), .B1 (n_878), .B2 (n_874));
OAI21_X1 i_673 (.ZN (n_5553), .A (n_859), .B1 (n_861), .B2 (n_857));
AOI21_X1 i_672 (.ZN (n_837), .A (n_5587), .B1 (n_5586), .B2 (n_843));
INV_X1 i_671 (.ZN (n_5590), .A (n_837));
AOI21_X1 i_670 (.ZN (n_5581), .A (n_888), .B1 (n_889), .B2 (n_886));
NAND2_X1 i_669 (.ZN (n_836), .A1 (inputB[20]), .A2 (inputA[27]));
INV_X1 i_668 (.ZN (n_835), .A (n_836));
NAND2_X1 i_667 (.ZN (n_834), .A1 (n_882), .A2 (n_835));
OAI21_X1 i_666 (.ZN (n_833), .A (n_834), .B1 (n_882), .B2 (n_835));
NAND2_X1 i_665 (.ZN (n_832), .A1 (inputB[22]), .A2 (inputA[25]));
XOR2_X1 i_664 (.Z (n_5660), .A (n_833), .B (n_832));
AOI22_X1 i_663 (.ZN (n_830), .A1 (inputB[24]), .A2 (inputA[23]), .B1 (inputB[23]), .B2 (inputA[24]));
INV_X1 i_662 (.ZN (n_829), .A (n_830));
NAND4_X1 i_661 (.ZN (n_828), .A1 (inputB[24]), .A2 (inputA[23]), .A3 (inputB[23]), .A4 (inputA[24]));
NAND2_X1 i_660 (.ZN (n_827), .A1 (n_829), .A2 (n_828));
NAND2_X1 i_659 (.ZN (n_826), .A1 (inputB[25]), .A2 (inputA[22]));
XOR2_X1 i_658 (.Z (n_5653), .A (n_827), .B (n_826));
NAND2_X1 i_657 (.ZN (n_825), .A1 (inputB[30]), .A2 (inputA[18]));
INV_X1 i_656 (.ZN (n_824), .A (n_825));
AOI22_X1 i_655 (.ZN (n_823), .A1 (inputB[30]), .A2 (inputA[17]), .B1 (inputB[29]), .B2 (inputA[18]));
AOI21_X1 i_654 (.ZN (n_822), .A (n_823), .B1 (n_872), .B2 (n_824));
NAND2_X1 i_653 (.ZN (n_821), .A1 (inputB[31]), .A2 (inputA[16]));
XOR2_X1 i_652 (.Z (n_5637), .A (n_822), .B (n_821));
AOI21_X1 i_651 (.ZN (n_820), .A (n_5592), .B1 (n_5591), .B2 (n_865));
INV_X1 i_650 (.ZN (n_5595), .A (n_820));
OAI21_X1 i_649 (.ZN (n_819), .A (n_881), .B1 (n_885), .B2 (n_879));
XOR2_X1 i_648 (.Z (n_5674), .A (n_5672), .B (n_819));
AOI21_X1 i_647 (.ZN (n_818), .A (n_5602), .B1 (n_5601), .B2 (n_856));
INV_X1 i_646 (.ZN (n_5605), .A (n_818));
OAI21_X1 i_645 (.ZN (n_817), .A (n_851), .B1 (n_5762), .B2 (n_5751));
INV_X1 i_644 (.ZN (n_816), .A (n_817));
NAND2_X1 i_643 (.ZN (n_815), .A1 (inputB[18]), .A2 (inputA[30]));
OR3_X1 i_642 (.ZN (n_814), .A1 (n_5762), .A2 (n_5750), .A3 (n_815));
NAND2_X1 i_641 (.ZN (n_813), .A1 (n_817), .A2 (n_814));
NAND2_X1 i_640 (.ZN (n_812), .A1 (inputB[19]), .A2 (inputA[28]));
XOR2_X1 i_639 (.Z (n_811), .A (n_813), .B (n_812));
XOR2_X1 i_638 (.Z (n_5684), .A (n_5682), .B (n_811));
AOI21_X1 i_637 (.ZN (n_810), .A (n_5607), .B1 (n_5606), .B2 (n_842));
INV_X1 i_636 (.ZN (n_5610), .A (n_810));
NAND2_X1 i_635 (.ZN (n_809), .A1 (inputB[28]), .A2 (inputA[19]));
AOI22_X1 i_634 (.ZN (n_808), .A1 (inputB[27]), .A2 (inputA[20]), .B1 (inputB[26]), .B2 (inputA[21]));
NAND2_X1 i_633 (.ZN (n_807), .A1 (inputB[27]), .A2 (inputA[21]));
INV_X1 i_632 (.ZN (n_806), .A (n_807));
NAND3_X1 i_631 (.ZN (n_805), .A1 (inputB[26]), .A2 (inputA[20]), .A3 (n_806));
INV_X1 i_630 (.ZN (n_804), .A (n_805));
NOR2_X1 i_629 (.ZN (n_803), .A1 (n_808), .A2 (n_804));
XNOR2_X1 i_628 (.ZN (n_802), .A (n_809), .B (n_803));
XOR2_X1 i_627 (.Z (n_5689), .A (n_5687), .B (n_802));
NAND2_X1 i_626 (.ZN (n_801), .A1 (n_871), .A2 (n_867));
XOR2_X1 i_625 (.Z (n_800), .A (n_5677), .B (n_801));
XOR2_X1 i_624 (.Z (n_5694), .A (n_5692), .B (n_800));
AOI21_X1 i_623 (.ZN (n_799), .A (n_5617), .B1 (n_5616), .B2 (n_844));
INV_X1 i_622 (.ZN (n_5620), .A (n_799));
AOI21_X1 i_621 (.ZN (n_798), .A (n_5612), .B1 (n_5611), .B2 (n_853));
INV_X1 i_620 (.ZN (n_797), .A (n_798));
XNOR2_X1 i_619 (.ZN (n_5704), .A (n_5702), .B (n_798));
AOI21_X1 i_618 (.ZN (n_796), .A (n_5597), .B1 (n_5596), .B2 (n_845));
INV_X1 i_617 (.ZN (n_795), .A (n_796));
XNOR2_X1 i_616 (.ZN (n_794), .A (n_5697), .B (n_796));
XOR2_X1 i_615 (.Z (n_5709), .A (n_5707), .B (n_794));
AOI21_X1 i_614 (.ZN (n_793), .A (n_5528), .B1 (n_5527), .B2 (n_898));
INV_X1 i_613 (.ZN (n_792), .A (n_793));
AOI21_X1 i_612 (.ZN (n_791), .A (n_5627), .B1 (n_5626), .B2 (n_792));
INV_X1 i_611 (.ZN (n_5630), .A (n_791));
OAI21_X1 i_610 (.ZN (n_5668), .A (n_814), .B1 (n_816), .B2 (n_812));
AOI22_X1 i_609 (.ZN (n_5661), .A1 (n_883), .A2 (n_836), .B1 (n_834), .B2 (n_832));
OAI21_X1 i_608 (.ZN (n_5647), .A (n_805), .B1 (n_809), .B2 (n_808));
AOI21_X1 i_607 (.ZN (n_790), .A (n_821), .B1 (n_872), .B2 (n_824));
NOR2_X1 i_606 (.ZN (n_5638), .A1 (n_823), .A2 (n_790));
AOI21_X1 i_605 (.ZN (n_789), .A (n_5673), .B1 (n_5672), .B2 (n_819));
INV_X1 i_604 (.ZN (n_5676), .A (n_789));
OAI211_X1 i_603 (.ZN (n_788), .A (inputB[19]), .B (inputA[29]), .C1 (n_5762), .C2 (n_5753));
AOI211_X1 i_602 (.ZN (n_787), .A (n_5762), .B (n_5753), .C1 (inputB[19]), .C2 (inputA[29]));
INV_X1 i_601 (.ZN (n_786), .A (n_787));
NAND2_X1 i_600 (.ZN (n_785), .A1 (n_788), .A2 (n_786));
XOR2_X1 i_599 (.Z (n_5752), .A (n_815), .B (n_785));
AOI22_X1 i_598 (.ZN (n_784), .A1 (inputB[24]), .A2 (inputA[24]), .B1 (inputB[23]), .B2 (inputA[25]));
INV_X1 i_597 (.ZN (n_783), .A (n_784));
NAND4_X1 i_596 (.ZN (n_782), .A1 (inputB[24]), .A2 (inputA[24]), .A3 (inputB[23]), .A4 (inputA[25]));
NAND2_X1 i_595 (.ZN (n_781), .A1 (n_783), .A2 (n_782));
NAND2_X1 i_594 (.ZN (n_780), .A1 (inputB[25]), .A2 (inputA[23]));
XOR2_X1 i_593 (.Z (n_5739), .A (n_781), .B (n_780));
NAND2_X1 i_592 (.ZN (n_779), .A1 (inputB[26]), .A2 (inputA[22]));
INV_X1 i_591 (.ZN (n_778), .A (n_779));
NAND2_X1 i_590 (.ZN (n_777), .A1 (n_806), .A2 (n_778));
NAND2_X1 i_589 (.ZN (n_776), .A1 (n_807), .A2 (n_779));
AND2_X1 i_588 (.ZN (n_775), .A1 (n_777), .A2 (n_776));
AND2_X1 i_587 (.ZN (n_774), .A1 (inputB[28]), .A2 (inputA[20]));
XOR2_X1 i_586 (.Z (n_5732), .A (n_775), .B (n_774));
AOI21_X1 i_585 (.ZN (n_773), .A (n_5678), .B1 (n_5677), .B2 (n_801));
INV_X1 i_584 (.ZN (n_772), .A (n_773));
XNOR2_X1 i_583 (.ZN (n_5766), .A (n_5764), .B (n_773));
OAI21_X1 i_582 (.ZN (n_771), .A (n_828), .B1 (n_830), .B2 (n_826));
XOR2_X1 i_581 (.Z (n_5761), .A (n_5759), .B (n_771));
AOI21_X1 i_580 (.ZN (n_770), .A (n_5683), .B1 (n_5682), .B2 (n_811));
INV_X1 i_579 (.ZN (n_5686), .A (n_770));
AOI21_X1 i_578 (.ZN (n_769), .A (n_5698), .B1 (n_5697), .B2 (n_795));
INV_X1 i_577 (.ZN (n_5701), .A (n_769));
NAND2_X1 i_576 (.ZN (n_768), .A1 (inputB[29]), .A2 (inputA[19]));
INV_X1 i_575 (.ZN (n_767), .A (n_768));
NAND2_X1 i_574 (.ZN (n_766), .A1 (n_824), .A2 (n_767));
NAND2_X1 i_573 (.ZN (n_765), .A1 (n_825), .A2 (n_768));
NAND2_X1 i_572 (.ZN (n_764), .A1 (n_766), .A2 (n_765));
NAND2_X1 i_571 (.ZN (n_763), .A1 (inputB[31]), .A2 (inputA[17]));
NAND2_X1 i_570 (.ZN (n_762), .A1 (n_765), .A2 (n_763));
XNOR2_X1 i_569 (.ZN (n_761), .A (n_764), .B (n_763));
XOR2_X1 i_568 (.Z (n_381), .A (n_2), .B (n_761));
AOI22_X1 i_567 (.ZN (n_760), .A1 (inputB[21]), .A2 (inputA[27]), .B1 (inputB[20]), .B2 (inputA[28]));
INV_X1 i_566 (.ZN (n_759), .A (n_760));
NAND3_X1 i_565 (.ZN (n_758), .A1 (inputB[21]), .A2 (inputA[28]), .A3 (n_835));
NAND2_X1 i_564 (.ZN (n_757), .A1 (n_759), .A2 (n_758));
NAND2_X1 i_563 (.ZN (n_756), .A1 (inputB[22]), .A2 (inputA[26]));
XOR2_X1 i_562 (.Z (n_755), .A (n_757), .B (n_756));
XOR2_X1 i_561 (.Z (n_380), .A (n_0), .B (n_755));
AOI21_X1 i_560 (.ZN (n_754), .A (n_5688), .B1 (n_5687), .B2 (n_802));
INV_X1 i_559 (.ZN (n_753), .A (n_754));
XNOR2_X1 i_558 (.ZN (n_379), .A (n_4), .B (n_754));
AOI21_X1 i_557 (.ZN (n_752), .A (n_5693), .B1 (n_5692), .B2 (n_800));
INV_X1 i_556 (.ZN (n_751), .A (n_752));
XNOR2_X1 i_555 (.ZN (n_378), .A (n_6), .B (n_752));
AOI21_X1 i_554 (.ZN (n_750), .A (n_5703), .B1 (n_5702), .B2 (n_797));
INV_X1 i_553 (.ZN (n_749), .A (n_750));
XNOR2_X1 i_552 (.ZN (n_377), .A (n_8), .B (n_750));
AOI21_X1 i_551 (.ZN (n_748), .A (n_5622), .B1 (n_5621), .B2 (n_841));
INV_X1 i_550 (.ZN (n_747), .A (n_748));
AOI21_X1 i_549 (.ZN (n_746), .A (n_5713), .B1 (n_5712), .B2 (n_747));
INV_X1 i_548 (.ZN (n_5716), .A (n_746));
OAI21_X1 i_547 (.ZN (n_5747), .A (n_758), .B1 (n_760), .B2 (n_756));
OAI21_X1 i_546 (.ZN (n_5740), .A (n_782), .B1 (n_784), .B2 (n_780));
NAND2_X1 i_545 (.ZN (n_5724), .A1 (n_766), .A2 (n_762));
AOI21_X1 i_544 (.ZN (n_745), .A (n_5760), .B1 (n_5759), .B2 (n_771));
INV_X1 i_543 (.ZN (n_5763), .A (n_745));
AOI22_X1 i_542 (.ZN (n_744), .A1 (inputB[21]), .A2 (inputA[28]), .B1 (inputB[20]), .B2 (inputA[29]));
INV_X1 i_541 (.ZN (n_743), .A (n_744));
NAND2_X1 i_540 (.ZN (n_742), .A1 (inputB[21]), .A2 (inputA[29]));
INV_X1 i_539 (.ZN (n_741), .A (n_742));
NAND3_X1 i_538 (.ZN (n_740), .A1 (inputB[20]), .A2 (inputA[28]), .A3 (n_741));
NAND2_X1 i_537 (.ZN (n_739), .A1 (n_743), .A2 (n_740));
NAND2_X1 i_536 (.ZN (n_738), .A1 (inputB[22]), .A2 (inputA[27]));
XOR2_X1 i_535 (.Z (n_376), .A (n_739), .B (n_738));
AND2_X1 i_534 (.ZN (n_737), .A1 (inputB[23]), .A2 (inputA[26]));
AOI21_X1 i_533 (.ZN (n_736), .A (n_737), .B1 (inputB[24]), .B2 (inputA[25]));
INV_X1 i_532 (.ZN (n_734), .A (n_736));
NAND3_X1 i_531 (.ZN (n_733), .A1 (inputB[24]), .A2 (inputA[25]), .A3 (n_737));
NAND2_X1 i_530 (.ZN (n_732), .A1 (n_734), .A2 (n_733));
NAND2_X1 i_529 (.ZN (n_731), .A1 (inputB[25]), .A2 (inputA[24]));
XOR2_X1 i_528 (.Z (n_375), .A (n_732), .B (n_731));
AOI22_X1 i_527 (.ZN (n_730), .A1 (inputB[30]), .A2 (inputA[19]), .B1 (inputB[29]), .B2 (inputA[20]));
INV_X1 i_526 (.ZN (n_729), .A (n_730));
NAND3_X1 i_525 (.ZN (n_728), .A1 (inputB[30]), .A2 (inputA[20]), .A3 (n_767));
NAND2_X1 i_524 (.ZN (n_727), .A1 (n_729), .A2 (n_728));
AND2_X1 i_523 (.ZN (n_726), .A1 (inputB[31]), .A2 (inputA[18]));
XOR2_X1 i_522 (.Z (n_374), .A (n_727), .B (n_726));
AOI21_X1 i_521 (.ZN (n_725), .A (n_5765), .B1 (n_5764), .B2 (n_772));
INV_X1 i_520 (.ZN (n_373), .A (n_725));
AOI21_X1 i_519 (.ZN (n_724), .A (n_3), .B1 (n_2), .B2 (n_761));
INV_X1 i_518 (.ZN (n_372), .A (n_724));
AOI21_X1 i_517 (.ZN (n_723), .A (n_1), .B1 (n_0), .B2 (n_755));
INV_X1 i_516 (.ZN (n_371), .A (n_723));
AOI21_X1 i_515 (.ZN (n_722), .A (n_5), .B1 (n_4), .B2 (n_753));
INV_X1 i_514 (.ZN (n_370), .A (n_722));
NAND2_X1 i_513 (.ZN (n_721), .A1 (inputB[27]), .A2 (inputA[23]));
INV_X1 i_512 (.ZN (n_720), .A (n_721));
NAND2_X1 i_511 (.ZN (n_719), .A1 (n_778), .A2 (n_720));
AOI22_X1 i_510 (.ZN (n_718), .A1 (inputB[27]), .A2 (inputA[22]), .B1 (inputB[26]), .B2 (inputA[23]));
INV_X1 i_509 (.ZN (n_717), .A (n_718));
NAND2_X1 i_508 (.ZN (n_716), .A1 (n_719), .A2 (n_717));
NAND2_X1 i_507 (.ZN (n_715), .A1 (inputB[28]), .A2 (inputA[21]));
XOR2_X1 i_506 (.Z (n_714), .A (n_716), .B (n_715));
XOR2_X1 i_505 (.Z (n_369), .A (n_18), .B (n_714));
AOI21_X1 i_504 (.ZN (n_713), .A (n_7), .B1 (n_6), .B2 (n_751));
INV_X1 i_503 (.ZN (n_368), .A (n_713));
NAND2_X1 i_502 (.ZN (n_712), .A1 (inputB[18]), .A2 (inputA[31]));
AND2_X1 i_501 (.ZN (n_711), .A1 (inputB[19]), .A2 (inputA[30]));
NAND2_X1 i_500 (.ZN (n_710), .A1 (n_712), .A2 (n_711));
OAI21_X1 i_499 (.ZN (n_709), .A (n_710), .B1 (n_712), .B2 (n_711));
AOI21_X1 i_498 (.ZN (n_708), .A (n_787), .B1 (n_815), .B2 (n_788));
INV_X1 i_497 (.ZN (n_707), .A (n_708));
XNOR2_X1 i_496 (.ZN (n_706), .A (n_709), .B (n_708));
XOR2_X1 i_495 (.Z (n_705), .A (n_16), .B (n_706));
XOR2_X1 i_494 (.Z (n_367), .A (n_22), .B (n_705));
NAND2_X1 i_493 (.ZN (n_704), .A1 (n_776), .A2 (n_774));
NAND2_X1 i_492 (.ZN (n_703), .A1 (n_777), .A2 (n_704));
XOR2_X1 i_491 (.Z (n_702), .A (n_14), .B (n_703));
XOR2_X1 i_490 (.Z (n_701), .A (n_20), .B (n_702));
XOR2_X1 i_489 (.Z (n_366), .A (n_24), .B (n_701));
AOI21_X1 i_488 (.ZN (n_700), .A (n_5708), .B1 (n_5707), .B2 (n_794));
INV_X1 i_487 (.ZN (n_699), .A (n_700));
AOI21_X1 i_486 (.ZN (n_698), .A (n_11), .B1 (n_10), .B2 (n_699));
INV_X1 i_485 (.ZN (n_365), .A (n_698));
NAND2_X1 i_484 (.ZN (n_639), .A1 (inputB[19]), .A2 (inputA[31]));
OAI21_X1 i_483 (.ZN (n_364), .A (n_740), .B1 (n_744), .B2 (n_738));
OAI21_X1 i_482 (.ZN (n_363), .A (n_719), .B1 (n_718), .B2 (n_715));
OAI21_X1 i_481 (.ZN (n_362), .A (n_728), .B1 (n_730), .B2 (n_726));
OAI21_X1 i_480 (.ZN (n_361), .A (n_710), .B1 (n_709), .B2 (n_707));
NAND3_X1 i_479 (.ZN (n_697), .A1 (inputB[20]), .A2 (inputA[30]), .A3 (n_741));
INV_X1 i_478 (.ZN (n_696), .A (n_697));
AOI21_X1 i_477 (.ZN (n_695), .A (n_741), .B1 (inputB[20]), .B2 (inputA[30]));
NOR2_X1 i_476 (.ZN (n_694), .A1 (n_696), .A2 (n_695));
NAND2_X1 i_475 (.ZN (n_693), .A1 (inputB[22]), .A2 (inputA[28]));
XNOR2_X1 i_474 (.ZN (n_360), .A (n_694), .B (n_693));
NAND2_X1 i_473 (.ZN (n_692), .A1 (inputB[26]), .A2 (inputA[24]));
INV_X1 i_472 (.ZN (n_691), .A (n_692));
NAND2_X1 i_471 (.ZN (n_690), .A1 (n_720), .A2 (n_691));
OAI21_X1 i_470 (.ZN (n_689), .A (n_690), .B1 (n_720), .B2 (n_691));
NAND2_X1 i_469 (.ZN (n_688), .A1 (inputB[28]), .A2 (inputA[22]));
XOR2_X1 i_468 (.Z (n_359), .A (n_689), .B (n_688));
AND2_X1 i_467 (.ZN (n_687), .A1 (inputB[31]), .A2 (inputA[19]));
AOI22_X1 i_466 (.ZN (n_686), .A1 (inputB[30]), .A2 (inputA[20]), .B1 (inputB[29]), .B2 (inputA[21]));
NAND2_X1 i_465 (.ZN (n_685), .A1 (inputB[30]), .A2 (inputA[21]));
INV_X1 i_464 (.ZN (n_684), .A (n_685));
NAND3_X1 i_463 (.ZN (n_683), .A1 (inputB[29]), .A2 (inputA[20]), .A3 (n_684));
INV_X1 i_462 (.ZN (n_682), .A (n_683));
NOR2_X1 i_461 (.ZN (n_681), .A1 (n_686), .A2 (n_682));
XNOR2_X1 i_460 (.ZN (n_358), .A (n_687), .B (n_681));
OAI21_X1 i_459 (.ZN (n_680), .A (n_733), .B1 (n_736), .B2 (n_731));
XOR2_X1 i_458 (.Z (n_357), .A (n_30), .B (n_680));
AOI21_X1 i_457 (.ZN (n_679), .A (n_19), .B1 (n_18), .B2 (n_714));
INV_X1 i_456 (.ZN (n_356), .A (n_679));
AOI21_X1 i_455 (.ZN (n_678), .A (n_21), .B1 (n_20), .B2 (n_702));
INV_X1 i_454 (.ZN (n_355), .A (n_678));
AOI21_X1 i_453 (.ZN (n_677), .A (n_15), .B1 (n_14), .B2 (n_703));
INV_X1 i_452 (.ZN (n_676), .A (n_677));
XNOR2_X1 i_451 (.ZN (n_675), .A (n_32), .B (n_677));
XOR2_X1 i_450 (.Z (n_354), .A (n_36), .B (n_675));
AOI21_X1 i_449 (.ZN (n_674), .A (n_23), .B1 (n_22), .B2 (n_705));
INV_X1 i_448 (.ZN (n_353), .A (n_674));
AOI21_X1 i_447 (.ZN (n_673), .A (n_17), .B1 (n_16), .B2 (n_706));
INV_X1 i_446 (.ZN (n_672), .A (n_673));
XNOR2_X1 i_445 (.ZN (n_352), .A (n_38), .B (n_673));
AOI21_X1 i_444 (.ZN (n_671), .A (n_9), .B1 (n_8), .B2 (n_749));
INV_X1 i_443 (.ZN (n_670), .A (n_671));
AOI21_X1 i_442 (.ZN (n_669), .A (n_27), .B1 (n_26), .B2 (n_670));
INV_X1 i_441 (.ZN (n_351), .A (n_669));
NAND2_X1 i_440 (.ZN (n_668), .A1 (inputB[24]), .A2 (inputA[27]));
INV_X1 i_439 (.ZN (n_667), .A (n_668));
NAND2_X1 i_438 (.ZN (n_666), .A1 (n_737), .A2 (n_667));
AOI22_X1 i_437 (.ZN (n_665), .A1 (inputB[24]), .A2 (inputA[26]), .B1 (inputB[23]), .B2 (inputA[27]));
INV_X1 i_436 (.ZN (n_664), .A (n_665));
NAND2_X1 i_435 (.ZN (n_663), .A1 (n_666), .A2 (n_664));
NAND2_X1 i_434 (.ZN (n_662), .A1 (inputB[25]), .A2 (inputA[25]));
XOR2_X1 i_433 (.Z (n_661), .A (n_663), .B (n_662));
XOR2_X1 i_432 (.Z (n_660), .A (n_34), .B (n_661));
XOR2_X1 i_431 (.Z (n_350), .A (n_40), .B (n_660));
OAI21_X1 i_430 (.ZN (n_349), .A (n_697), .B1 (n_695), .B2 (n_693));
OAI21_X1 i_429 (.ZN (n_348), .A (n_666), .B1 (n_665), .B2 (n_662));
AOI21_X1 i_428 (.ZN (n_347), .A (n_686), .B1 (n_687), .B2 (n_683));
AOI21_X1 i_427 (.ZN (n_659), .A (n_31), .B1 (n_30), .B2 (n_680));
INV_X1 i_426 (.ZN (n_346), .A (n_659));
NAND2_X1 i_425 (.ZN (n_658), .A1 (inputB[23]), .A2 (inputA[28]));
INV_X1 i_424 (.ZN (n_657), .A (n_658));
NAND2_X1 i_423 (.ZN (n_656), .A1 (n_667), .A2 (n_657));
NAND2_X1 i_422 (.ZN (n_655), .A1 (n_668), .A2 (n_658));
AND2_X1 i_421 (.ZN (n_654), .A1 (n_656), .A2 (n_655));
AND2_X1 i_420 (.ZN (n_653), .A1 (inputB[25]), .A2 (inputA[26]));
XOR2_X1 i_419 (.Z (n_345), .A (n_654), .B (n_653));
AOI22_X1 i_418 (.ZN (n_652), .A1 (inputB[27]), .A2 (inputA[24]), .B1 (inputB[26]), .B2 (inputA[25]));
INV_X1 i_417 (.ZN (n_651), .A (n_652));
NAND3_X1 i_416 (.ZN (n_650), .A1 (inputB[27]), .A2 (inputA[25]), .A3 (n_691));
NAND2_X1 i_415 (.ZN (n_649), .A1 (n_651), .A2 (n_650));
NAND2_X1 i_414 (.ZN (n_648), .A1 (inputB[28]), .A2 (inputA[23]));
XOR2_X1 i_413 (.Z (n_344), .A (n_649), .B (n_648));
AOI21_X1 i_412 (.ZN (n_647), .A (n_33), .B1 (n_32), .B2 (n_676));
INV_X1 i_411 (.ZN (n_343), .A (n_647));
AOI22_X1 i_410 (.ZN (n_646), .A1 (n_721), .A2 (n_692), .B1 (n_690), .B2 (n_688));
XOR2_X1 i_409 (.Z (n_342), .A (n_46), .B (n_646));
NAND2_X1 i_408 (.ZN (n_645), .A1 (inputB[22]), .A2 (inputA[30]));
NOR2_X1 i_407 (.ZN (n_644), .A1 (n_742), .A2 (n_645));
AOI22_X1 i_406 (.ZN (n_643), .A1 (inputB[21]), .A2 (inputA[30]), .B1 (inputB[22]), .B2 (inputA[29]));
INV_X1 i_405 (.ZN (n_642), .A (n_643));
NOR2_X1 i_404 (.ZN (n_641), .A1 (n_644), .A2 (n_643));
NAND2_X1 i_403 (.ZN (n_640), .A1 (inputB[20]), .A2 (inputA[31]));
XOR2_X1 i_402 (.Z (n_638), .A (n_641), .B (n_640));
XOR2_X1 i_401 (.Z (n_341), .A (n_48), .B (n_638));
AOI21_X1 i_400 (.ZN (n_637), .A (n_39), .B1 (n_38), .B2 (n_672));
INV_X1 i_399 (.ZN (n_340), .A (n_637));
NAND2_X1 i_398 (.ZN (n_636), .A1 (inputB[29]), .A2 (inputA[22]));
INV_X1 i_397 (.ZN (n_635), .A (n_636));
NAND2_X1 i_396 (.ZN (n_634), .A1 (n_684), .A2 (n_635));
NAND2_X1 i_395 (.ZN (n_633), .A1 (n_685), .A2 (n_636));
NAND2_X1 i_394 (.ZN (n_632), .A1 (n_634), .A2 (n_633));
NAND2_X1 i_393 (.ZN (n_631), .A1 (inputB[31]), .A2 (inputA[20]));
NAND2_X1 i_392 (.ZN (n_630), .A1 (n_633), .A2 (n_631));
XNOR2_X1 i_391 (.ZN (n_629), .A (n_632), .B (n_631));
XOR2_X1 i_390 (.Z (n_339), .A (n_50), .B (n_629));
AOI21_X1 i_389 (.ZN (n_628), .A (n_35), .B1 (n_34), .B2 (n_661));
INV_X1 i_388 (.ZN (n_627), .A (n_628));
XNOR2_X1 i_387 (.ZN (n_338), .A (n_52), .B (n_628));
AOI21_X1 i_386 (.ZN (n_626), .A (n_37), .B1 (n_36), .B2 (n_675));
INV_X1 i_385 (.ZN (n_625), .A (n_626));
XNOR2_X1 i_384 (.ZN (n_337), .A (n_54), .B (n_626));
AOI21_X1 i_383 (.ZN (n_624), .A (n_25), .B1 (n_24), .B2 (n_701));
INV_X1 i_382 (.ZN (n_623), .A (n_624));
AOI21_X1 i_381 (.ZN (n_622), .A (n_43), .B1 (n_42), .B2 (n_623));
INV_X1 i_380 (.ZN (n_336), .A (n_622));
NAND2_X1 i_379 (.ZN (n_621), .A1 (n_655), .A2 (n_653));
NAND2_X1 i_378 (.ZN (n_335), .A1 (n_656), .A2 (n_621));
OAI21_X1 i_377 (.ZN (n_334), .A (n_650), .B1 (n_652), .B2 (n_648));
AOI21_X1 i_376 (.ZN (n_620), .A (n_47), .B1 (n_46), .B2 (n_646));
INV_X1 i_375 (.ZN (n_333), .A (n_620));
AOI21_X1 i_374 (.ZN (n_619), .A (n_644), .B1 (n_642), .B2 (n_640));
INV_X1 i_373 (.ZN (n_618), .A (n_619));
NAND2_X1 i_372 (.ZN (n_617), .A1 (inputB[21]), .A2 (inputA[31]));
XNOR2_X1 i_371 (.ZN (n_616), .A (n_645), .B (n_617));
XOR2_X1 i_370 (.Z (n_332), .A (n_618), .B (n_616));
AOI22_X1 i_369 (.ZN (n_615), .A1 (inputB[27]), .A2 (inputA[25]), .B1 (inputB[26]), .B2 (inputA[26]));
INV_X1 i_368 (.ZN (n_614), .A (n_615));
NAND2_X1 i_367 (.ZN (n_613), .A1 (inputB[27]), .A2 (inputA[26]));
INV_X1 i_366 (.ZN (n_612), .A (n_613));
NAND3_X1 i_365 (.ZN (n_611), .A1 (inputB[26]), .A2 (inputA[25]), .A3 (n_612));
NAND2_X1 i_364 (.ZN (n_610), .A1 (n_614), .A2 (n_611));
NAND2_X1 i_363 (.ZN (n_609), .A1 (inputB[28]), .A2 (inputA[24]));
XOR2_X1 i_362 (.Z (n_331), .A (n_610), .B (n_609));
NAND2_X1 i_361 (.ZN (n_608), .A1 (inputB[30]), .A2 (inputA[23]));
INV_X1 i_360 (.ZN (n_607), .A (n_608));
AOI22_X1 i_359 (.ZN (n_606), .A1 (inputB[30]), .A2 (inputA[22]), .B1 (inputB[29]), .B2 (inputA[23]));
AOI21_X1 i_358 (.ZN (n_605), .A (n_606), .B1 (n_635), .B2 (n_607));
NAND2_X1 i_357 (.ZN (n_604), .A1 (inputB[31]), .A2 (inputA[21]));
XOR2_X1 i_356 (.Z (n_330), .A (n_605), .B (n_604));
AOI21_X1 i_355 (.ZN (n_603), .A (n_51), .B1 (n_50), .B2 (n_629));
INV_X1 i_354 (.ZN (n_329), .A (n_603));
AOI21_X1 i_353 (.ZN (n_602), .A (n_49), .B1 (n_48), .B2 (n_638));
INV_X1 i_352 (.ZN (n_328), .A (n_602));
NAND2_X1 i_351 (.ZN (n_601), .A1 (n_634), .A2 (n_630));
XOR2_X1 i_350 (.Z (n_600), .A (n_60), .B (n_601));
XOR2_X1 i_349 (.Z (n_327), .A (n_64), .B (n_600));
NOR2_X1 i_348 (.ZN (n_599), .A1 (n_5767), .A2 (n_5750));
NAND2_X1 i_347 (.ZN (n_598), .A1 (n_657), .A2 (n_599));
AOI22_X1 i_346 (.ZN (n_597), .A1 (inputB[24]), .A2 (inputA[28]), .B1 (inputB[23]), .B2 (inputA[29]));
INV_X1 i_345 (.ZN (n_596), .A (n_597));
NAND2_X1 i_344 (.ZN (n_595), .A1 (n_598), .A2 (n_596));
NAND2_X1 i_343 (.ZN (n_594), .A1 (inputB[25]), .A2 (inputA[27]));
XOR2_X1 i_342 (.Z (n_593), .A (n_595), .B (n_594));
XOR2_X1 i_341 (.Z (n_326), .A (n_62), .B (n_593));
AOI21_X1 i_340 (.ZN (n_592), .A (n_53), .B1 (n_52), .B2 (n_627));
INV_X1 i_339 (.ZN (n_591), .A (n_592));
XNOR2_X1 i_338 (.ZN (n_325), .A (n_66), .B (n_592));
AOI21_X1 i_337 (.ZN (n_590), .A (n_41), .B1 (n_40), .B2 (n_660));
INV_X1 i_336 (.ZN (n_589), .A (n_590));
AOI21_X1 i_335 (.ZN (n_588), .A (n_57), .B1 (n_56), .B2 (n_589));
INV_X1 i_334 (.ZN (n_324), .A (n_588));
NAND2_X1 i_333 (.ZN (n_735), .A1 (inputB[22]), .A2 (inputA[31]));
OAI21_X1 i_332 (.ZN (n_323), .A (n_598), .B1 (n_597), .B2 (n_594));
AOI21_X1 i_331 (.ZN (n_587), .A (n_604), .B1 (n_635), .B2 (n_607));
NOR2_X1 i_330 (.ZN (n_322), .A1 (n_606), .A2 (n_587));
AOI21_X1 i_329 (.ZN (n_586), .A (n_61), .B1 (n_60), .B2 (n_601));
INV_X1 i_328 (.ZN (n_321), .A (n_586));
AOI21_X1 i_327 (.ZN (n_585), .A (n_599), .B1 (inputB[23]), .B2 (inputA[30]));
INV_X1 i_326 (.ZN (n_584), .A (n_585));
NAND3_X1 i_325 (.ZN (n_583), .A1 (inputB[23]), .A2 (inputA[30]), .A3 (n_599));
NAND2_X1 i_324 (.ZN (n_582), .A1 (n_584), .A2 (n_583));
NAND2_X1 i_323 (.ZN (n_581), .A1 (inputB[25]), .A2 (inputA[28]));
XOR2_X1 i_322 (.Z (n_320), .A (n_582), .B (n_581));
NAND2_X1 i_321 (.ZN (n_580), .A1 (inputB[26]), .A2 (inputA[27]));
INV_X1 i_320 (.ZN (n_579), .A (n_580));
NAND2_X1 i_319 (.ZN (n_578), .A1 (n_612), .A2 (n_579));
OAI21_X1 i_318 (.ZN (n_577), .A (n_578), .B1 (n_612), .B2 (n_579));
NAND2_X1 i_317 (.ZN (n_576), .A1 (inputB[28]), .A2 (inputA[25]));
XOR2_X1 i_316 (.Z (n_319), .A (n_577), .B (n_576));
OAI21_X1 i_315 (.ZN (n_575), .A (n_611), .B1 (n_615), .B2 (n_609));
XOR2_X1 i_314 (.Z (n_318), .A (n_72), .B (n_575));
AOI21_X1 i_313 (.ZN (n_574), .A (n_63), .B1 (n_62), .B2 (n_593));
INV_X1 i_312 (.ZN (n_317), .A (n_574));
AOI21_X1 i_311 (.ZN (n_573), .A (n_65), .B1 (n_64), .B2 (n_600));
INV_X1 i_310 (.ZN (n_316), .A (n_573));
NAND2_X1 i_309 (.ZN (n_572), .A1 (inputB[29]), .A2 (inputA[24]));
INV_X1 i_308 (.ZN (n_571), .A (n_572));
NAND2_X1 i_307 (.ZN (n_570), .A1 (n_607), .A2 (n_571));
NAND2_X1 i_306 (.ZN (n_569), .A1 (n_608), .A2 (n_572));
AND2_X1 i_305 (.ZN (n_568), .A1 (n_570), .A2 (n_569));
NAND2_X1 i_304 (.ZN (n_567), .A1 (inputB[31]), .A2 (inputA[22]));
XOR2_X1 i_303 (.Z (n_566), .A (n_568), .B (n_567));
XOR2_X1 i_302 (.Z (n_315), .A (n_76), .B (n_566));
AOI21_X1 i_301 (.ZN (n_565), .A (n_645), .B1 (n_619), .B2 (n_616));
AOI21_X1 i_300 (.ZN (n_564), .A (n_565), .B1 (n_618), .B2 (n_617));
INV_X1 i_299 (.ZN (n_563), .A (n_564));
XNOR2_X1 i_298 (.ZN (n_562), .A (n_74), .B (n_564));
XOR2_X1 i_297 (.Z (n_314), .A (n_78), .B (n_562));
AOI21_X1 i_296 (.ZN (n_561), .A (n_55), .B1 (n_54), .B2 (n_625));
INV_X1 i_295 (.ZN (n_560), .A (n_561));
AOI21_X1 i_294 (.ZN (n_559), .A (n_69), .B1 (n_68), .B2 (n_560));
INV_X1 i_293 (.ZN (n_313), .A (n_559));
OAI21_X1 i_292 (.ZN (n_312), .A (n_583), .B1 (n_585), .B2 (n_581));
AOI22_X1 i_291 (.ZN (n_311), .A1 (n_613), .A2 (n_580), .B1 (n_578), .B2 (n_576));
AOI21_X1 i_290 (.ZN (n_558), .A (n_73), .B1 (n_72), .B2 (n_575));
INV_X1 i_289 (.ZN (n_310), .A (n_558));
NAND2_X1 i_288 (.ZN (n_557), .A1 (inputB[23]), .A2 (inputA[31]));
NAND3_X1 i_287 (.ZN (n_556), .A1 (inputB[24]), .A2 (inputA[30]), .A3 (n_557));
INV_X1 i_286 (.ZN (n_555), .A (n_556));
AOI21_X1 i_285 (.ZN (n_554), .A (n_557), .B1 (inputB[24]), .B2 (inputA[30]));
NOR2_X1 i_284 (.ZN (n_553), .A1 (n_555), .A2 (n_554));
NAND2_X1 i_283 (.ZN (n_552), .A1 (inputB[25]), .A2 (inputA[29]));
XNOR2_X1 i_282 (.ZN (n_309), .A (n_553), .B (n_552));
AND2_X1 i_281 (.ZN (n_551), .A1 (inputB[30]), .A2 (inputA[25]));
AOI22_X1 i_280 (.ZN (n_550), .A1 (inputB[30]), .A2 (inputA[24]), .B1 (inputB[29]), .B2 (inputA[25]));
AOI21_X1 i_279 (.ZN (n_549), .A (n_550), .B1 (n_571), .B2 (n_551));
NAND2_X1 i_278 (.ZN (n_548), .A1 (inputB[31]), .A2 (inputA[23]));
XOR2_X1 i_277 (.Z (n_308), .A (n_549), .B (n_548));
AOI21_X1 i_276 (.ZN (n_547), .A (n_75), .B1 (n_74), .B2 (n_563));
INV_X1 i_275 (.ZN (n_307), .A (n_547));
AOI21_X1 i_274 (.ZN (n_546), .A (n_77), .B1 (n_76), .B2 (n_566));
INV_X1 i_273 (.ZN (n_306), .A (n_546));
NAND2_X1 i_272 (.ZN (n_545), .A1 (inputB[27]), .A2 (inputA[28]));
INV_X1 i_271 (.ZN (n_544), .A (n_545));
NAND2_X1 i_270 (.ZN (n_542), .A1 (n_579), .A2 (n_544));
AOI22_X1 i_269 (.ZN (n_541), .A1 (inputB[27]), .A2 (inputA[27]), .B1 (inputB[26]), .B2 (inputA[28]));
INV_X1 i_268 (.ZN (n_540), .A (n_541));
NAND2_X1 i_267 (.ZN (n_539), .A1 (n_542), .A2 (n_540));
NAND2_X1 i_266 (.ZN (n_538), .A1 (inputB[28]), .A2 (inputA[26]));
XOR2_X1 i_265 (.Z (n_537), .A (n_539), .B (n_538));
XOR2_X1 i_264 (.Z (n_305), .A (n_86), .B (n_537));
AOI21_X1 i_263 (.ZN (n_536), .A (n_79), .B1 (n_78), .B2 (n_562));
INV_X1 i_262 (.ZN (n_304), .A (n_536));
AOI21_X1 i_261 (.ZN (n_535), .A (n_67), .B1 (n_66), .B2 (n_591));
INV_X1 i_260 (.ZN (n_534), .A (n_535));
AOI21_X1 i_259 (.ZN (n_533), .A (n_81), .B1 (n_80), .B2 (n_534));
INV_X1 i_258 (.ZN (n_303), .A (n_533));
OAI21_X1 i_257 (.ZN (n_302), .A (n_542), .B1 (n_541), .B2 (n_538));
AOI22_X1 i_256 (.ZN (n_532), .A1 (n_571), .A2 (n_551), .B1 (n_549), .B2 (n_548));
INV_X1 i_255 (.ZN (n_301), .A (n_532));
AOI211_X1 i_254 (.ZN (n_531), .A (n_5767), .B (n_5753), .C1 (inputB[25]), .C2 (inputA[30]));
OAI211_X1 i_253 (.ZN (n_530), .A (inputB[25]), .B (inputA[30]), .C1 (n_5767), .C2 (n_5753));
INV_X1 i_252 (.ZN (n_529), .A (n_530));
NOR2_X1 i_251 (.ZN (n_528), .A1 (n_531), .A2 (n_529));
AOI21_X1 i_250 (.ZN (n_527), .A (n_554), .B1 (n_556), .B2 (n_552));
INV_X1 i_249 (.ZN (n_526), .A (n_527));
XOR2_X1 i_248 (.Z (n_300), .A (n_528), .B (n_527));
NAND2_X1 i_247 (.ZN (n_525), .A1 (inputB[26]), .A2 (inputA[29]));
INV_X1 i_246 (.ZN (n_524), .A (n_525));
NAND2_X1 i_245 (.ZN (n_523), .A1 (n_544), .A2 (n_524));
OAI21_X1 i_244 (.ZN (n_522), .A (n_523), .B1 (n_544), .B2 (n_524));
NAND2_X1 i_243 (.ZN (n_521), .A1 (inputB[28]), .A2 (inputA[27]));
XOR2_X1 i_242 (.Z (n_299), .A (n_522), .B (n_521));
NAND2_X1 i_241 (.ZN (n_520), .A1 (n_569), .A2 (n_567));
NAND2_X1 i_240 (.ZN (n_519), .A1 (n_570), .A2 (n_520));
AOI21_X1 i_239 (.ZN (n_518), .A (n_85), .B1 (n_84), .B2 (n_519));
INV_X1 i_238 (.ZN (n_517), .A (n_518));
XNOR2_X1 i_237 (.ZN (n_298), .A (n_94), .B (n_518));
AOI21_X1 i_236 (.ZN (n_516), .A (n_87), .B1 (n_86), .B2 (n_537));
INV_X1 i_235 (.ZN (n_297), .A (n_516));
AOI21_X1 i_234 (.ZN (n_515), .A (n_551), .B1 (inputB[29]), .B2 (inputA[26]));
NAND3_X1 i_233 (.ZN (n_514), .A1 (inputB[29]), .A2 (inputA[26]), .A3 (n_551));
INV_X1 i_232 (.ZN (n_513), .A (n_514));
NOR2_X1 i_231 (.ZN (n_512), .A1 (n_515), .A2 (n_513));
NAND2_X1 i_230 (.ZN (n_511), .A1 (inputB[31]), .A2 (inputA[24]));
INV_X1 i_229 (.ZN (n_510), .A (n_511));
XOR2_X1 i_228 (.Z (n_509), .A (n_512), .B (n_511));
XOR2_X1 i_227 (.Z (n_296), .A (n_96), .B (n_509));
XOR2_X1 i_226 (.Z (n_508), .A (n_84), .B (n_519));
AOI21_X1 i_225 (.ZN (n_507), .A (n_89), .B1 (n_88), .B2 (n_508));
INV_X1 i_224 (.ZN (n_506), .A (n_507));
XNOR2_X1 i_223 (.ZN (n_295), .A (n_98), .B (n_507));
NAND2_X1 i_222 (.ZN (n_831), .A1 (inputB[25]), .A2 (inputA[31]));
AOI22_X1 i_221 (.ZN (n_294), .A1 (n_545), .A2 (n_525), .B1 (n_523), .B2 (n_521));
AOI21_X1 i_220 (.ZN (n_293), .A (n_531), .B1 (n_530), .B2 (n_526));
AOI22_X1 i_219 (.ZN (n_505), .A1 (inputB[27]), .A2 (inputA[29]), .B1 (inputB[26]), .B2 (inputA[30]));
INV_X1 i_218 (.ZN (n_504), .A (n_505));
NAND2_X1 i_217 (.ZN (n_503), .A1 (inputB[27]), .A2 (inputA[30]));
OAI21_X1 i_216 (.ZN (n_502), .A (n_504), .B1 (n_525), .B2 (n_503));
NAND2_X1 i_215 (.ZN (n_501), .A1 (inputB[28]), .A2 (inputA[28]));
XOR2_X1 i_214 (.Z (n_292), .A (n_502), .B (n_501));
AOI21_X1 i_213 (.ZN (n_500), .A (n_95), .B1 (n_94), .B2 (n_517));
INV_X1 i_212 (.ZN (n_291), .A (n_500));
OAI21_X1 i_211 (.ZN (n_499), .A (n_514), .B1 (n_515), .B2 (n_510));
XOR2_X1 i_210 (.Z (n_290), .A (n_102), .B (n_499));
AND2_X1 i_209 (.ZN (n_498), .A1 (inputB[29]), .A2 (inputA[27]));
AOI21_X1 i_208 (.ZN (n_497), .A (n_498), .B1 (inputB[30]), .B2 (inputA[26]));
NAND3_X1 i_207 (.ZN (n_496), .A1 (inputB[30]), .A2 (inputA[26]), .A3 (n_498));
INV_X1 i_206 (.ZN (n_495), .A (n_496));
NOR2_X1 i_205 (.ZN (n_494), .A1 (n_497), .A2 (n_495));
AND2_X1 i_204 (.ZN (n_493), .A1 (inputB[31]), .A2 (inputA[25]));
XNOR2_X1 i_203 (.ZN (n_492), .A (n_494), .B (n_493));
XOR2_X1 i_202 (.Z (n_289), .A (n_104), .B (n_492));
AOI21_X1 i_201 (.ZN (n_491), .A (n_99), .B1 (n_98), .B2 (n_506));
INV_X1 i_200 (.ZN (n_288), .A (n_491));
OAI22_X1 i_199 (.ZN (n_287), .A1 (n_525), .A2 (n_503), .B1 (n_505), .B2 (n_501));
AOI21_X1 i_198 (.ZN (n_286), .A (n_497), .B1 (n_496), .B2 (n_493));
AOI21_X1 i_197 (.ZN (n_490), .A (n_503), .B1 (inputB[26]), .B2 (inputA[31]));
INV_X1 i_196 (.ZN (n_489), .A (n_490));
AND3_X1 i_195 (.ZN (n_488), .A1 (inputB[26]), .A2 (inputA[31]), .A3 (n_503));
NOR2_X1 i_194 (.ZN (n_487), .A1 (n_490), .A2 (n_488));
NAND2_X1 i_193 (.ZN (n_486), .A1 (inputB[28]), .A2 (inputA[29]));
XNOR2_X1 i_192 (.ZN (n_285), .A (n_487), .B (n_486));
NAND2_X1 i_191 (.ZN (n_485), .A1 (inputB[30]), .A2 (inputA[28]));
INV_X1 i_190 (.ZN (n_484), .A (n_485));
NAND2_X1 i_189 (.ZN (n_483), .A1 (n_498), .A2 (n_484));
AOI22_X1 i_188 (.ZN (n_482), .A1 (inputB[30]), .A2 (inputA[27]), .B1 (inputB[29]), .B2 (inputA[28]));
INV_X1 i_187 (.ZN (n_481), .A (n_482));
NAND2_X1 i_186 (.ZN (n_480), .A1 (n_483), .A2 (n_481));
NAND2_X1 i_185 (.ZN (n_479), .A1 (inputB[31]), .A2 (inputA[26]));
INV_X1 i_184 (.ZN (n_478), .A (n_479));
XNOR2_X1 i_183 (.ZN (n_284), .A (n_480), .B (n_479));
AOI21_X1 i_182 (.ZN (n_477), .A (n_105), .B1 (n_104), .B2 (n_492));
INV_X1 i_181 (.ZN (n_283), .A (n_477));
AOI21_X1 i_180 (.ZN (n_476), .A (n_97), .B1 (n_96), .B2 (n_509));
INV_X1 i_179 (.ZN (n_475), .A (n_476));
AOI21_X1 i_178 (.ZN (n_474), .A (n_107), .B1 (n_106), .B2 (n_475));
INV_X1 i_177 (.ZN (n_282), .A (n_474));
AOI21_X1 i_176 (.ZN (n_281), .A (n_482), .B1 (n_483), .B2 (n_478));
AOI21_X1 i_175 (.ZN (n_473), .A (n_488), .B1 (n_489), .B2 (n_486));
INV_X1 i_174 (.ZN (n_472), .A (n_473));
NAND2_X1 i_173 (.ZN (n_471), .A1 (inputB[28]), .A2 (inputA[30]));
NAND2_X1 i_172 (.ZN (n_470), .A1 (inputB[27]), .A2 (inputA[31]));
XNOR2_X1 i_171 (.ZN (n_469), .A (n_471), .B (n_470));
XOR2_X1 i_170 (.Z (n_280), .A (n_473), .B (n_469));
AOI21_X1 i_169 (.ZN (n_468), .A (n_103), .B1 (n_102), .B2 (n_499));
INV_X1 i_168 (.ZN (n_467), .A (n_468));
AOI21_X1 i_167 (.ZN (n_466), .A (n_111), .B1 (n_110), .B2 (n_467));
INV_X1 i_166 (.ZN (n_279), .A (n_466));
XNOR2_X1 i_165 (.ZN (n_465), .A (n_110), .B (n_468));
AOI21_X1 i_164 (.ZN (n_464), .A (n_113), .B1 (n_112), .B2 (n_465));
INV_X1 i_163 (.ZN (n_278), .A (n_464));
NAND2_X1 i_162 (.ZN (n_927), .A1 (inputB[28]), .A2 (inputA[31]));
NAND2_X1 i_161 (.ZN (n_463), .A1 (inputB[29]), .A2 (inputA[29]));
INV_X1 i_160 (.ZN (n_462), .A (n_463));
NAND2_X1 i_159 (.ZN (n_461), .A1 (n_484), .A2 (n_462));
AND2_X1 i_158 (.ZN (n_460), .A1 (inputB[31]), .A2 (inputA[27]));
AOI22_X1 i_157 (.ZN (n_277), .A1 (n_485), .A2 (n_463), .B1 (n_461), .B2 (n_460));
AOI22_X1 i_156 (.ZN (n_459), .A1 (inputB[30]), .A2 (inputA[29]), .B1 (inputB[29]), .B2 (inputA[30]));
AOI21_X1 i_155 (.ZN (n_458), .A (n_459), .B1 (n_5748), .B2 (n_462));
NAND2_X1 i_154 (.ZN (n_457), .A1 (inputB[31]), .A2 (inputA[28]));
XOR2_X1 i_153 (.Z (n_276), .A (n_458), .B (n_457));
AOI21_X1 i_152 (.ZN (n_456), .A (n_471), .B1 (n_472), .B2 (n_469));
AOI21_X1 i_151 (.ZN (n_455), .A (n_456), .B1 (n_473), .B2 (n_470));
INV_X1 i_150 (.ZN (n_454), .A (n_455));
XNOR2_X1 i_149 (.ZN (n_275), .A (n_120), .B (n_455));
AOI22_X1 i_148 (.ZN (n_453), .A1 (n_5748), .A2 (n_462), .B1 (n_458), .B2 (n_457));
INV_X1 i_147 (.ZN (n_274), .A (n_453));
XOR2_X1 i_146 (.Z (n_273), .A (n_5745), .B (n_5743));
NAND2_X1 i_145 (.ZN (n_1022), .A1 (inputB[31]), .A2 (inputA[30]));
NAND2_X1 i_144 (.ZN (n_991), .A1 (inputB[30]), .A2 (inputA[31]));
OAI22_X1 i_143 (.ZN (n_1034), .A1 (n_5495), .A2 (n_5477), .B1 (n_5496), .B2 (n_5478));
NAND2_X1 i_142 (.ZN (n_452), .A1 (n_5483), .A2 (n_5481));
XOR2_X1 i_141 (.Z (n_1029), .A (n_5480), .B (n_452));
NAND2_X1 i_140 (.ZN (n_451), .A1 (n_5470), .A2 (n_5466));
XOR2_X1 i_139 (.Z (n_1039), .A (n_5465), .B (n_451));
XOR2_X1 i_138 (.Z (n_1070), .A (n_1068), .B (n_5426));
XOR2_X1 i_137 (.Z (n_1099), .A (n_1097), .B (n_5368));
XOR2_X1 i_136 (.Z (n_1133), .A (n_1103), .B (n_1131));
XOR2_X1 i_135 (.Z (n_1171), .A (n_1137), .B (n_1169));
XOR2_X1 i_134 (.Z (n_1217), .A (n_1215), .B (n_5238));
XOR2_X1 i_133 (.Z (n_1268), .A (n_1266), .B (n_5159));
XOR2_X1 i_132 (.Z (n_1323), .A (n_1321), .B (n_5118));
XOR2_X1 i_131 (.Z (n_1386), .A (n_1384), .B (n_4956));
XNOR2_X1 i_130 (.ZN (n_1454), .A (n_1452), .B (n_4951));
XOR2_X1 i_129 (.Z (n_1526), .A (n_1524), .B (n_4873));
XOR2_X1 i_128 (.Z (n_1606), .A (n_1604), .B (n_4762));
XOR2_X1 i_127 (.Z (n_1691), .A (n_1689), .B (n_4655));
XOR2_X1 i_126 (.Z (n_1780), .A (n_1778), .B (n_4563));
XOR2_X1 i_125 (.Z (n_2085), .A (n_2083), .B (n_4205));
XOR2_X1 i_124 (.Z (n_2708), .A (n_2706), .B (n_3509));
AOI21_X1 i_123 (.ZN (n_450), .A (n_3641), .B1 (n_3640), .B2 (n_2644));
INV_X1 i_122 (.ZN (n_449), .A (n_450));
XNOR2_X1 i_121 (.ZN (n_3814), .A (n_3812), .B (n_450));
AOI21_X1 i_120 (.ZN (n_448), .A (n_3813), .B1 (n_3812), .B2 (n_449));
INV_X1 i_119 (.ZN (n_3816), .A (n_448));
XNOR2_X1 i_118 (.ZN (n_446), .A (n_3974), .B (n_2155));
XOR2_X1 i_117 (.Z (n_3981), .A (n_3979), .B (n_446));
AOI21_X1 i_116 (.ZN (n_445), .A (n_3980), .B1 (n_3979), .B2 (n_446));
INV_X1 i_115 (.ZN (n_3983), .A (n_445));
XNOR2_X1 i_114 (.ZN (n_444), .A (n_4136), .B (n_2018));
XOR2_X1 i_113 (.Z (n_4143), .A (n_4141), .B (n_444));
XOR2_X1 i_112 (.Z (n_443), .A (n_4290), .B (n_1868));
XOR2_X1 i_111 (.Z (n_4297), .A (n_4295), .B (n_443));
AOI21_X1 i_110 (.ZN (n_442), .A (n_4142), .B1 (n_4141), .B2 (n_444));
INV_X1 i_109 (.ZN (n_4145), .A (n_442));
AOI21_X1 i_108 (.ZN (n_441), .A (n_4296), .B1 (n_4295), .B2 (n_443));
INV_X1 i_107 (.ZN (n_4299), .A (n_441));
XNOR2_X1 i_106 (.ZN (n_440), .A (n_4440), .B (n_1725));
XOR2_X1 i_105 (.Z (n_4447), .A (n_4445), .B (n_440));
AOI21_X1 i_104 (.ZN (n_439), .A (n_4446), .B1 (n_4445), .B2 (n_440));
INV_X1 i_103 (.ZN (n_4449), .A (n_439));
XNOR2_X1 i_102 (.ZN (n_438), .A (n_4585), .B (n_1592));
XOR2_X1 i_101 (.Z (n_4592), .A (n_4590), .B (n_438));
AOI21_X1 i_100 (.ZN (n_437), .A (n_4591), .B1 (n_4590), .B2 (n_438));
INV_X1 i_99 (.ZN (n_4594), .A (n_437));
XNOR2_X1 i_98 (.ZN (n_436), .A (n_4722), .B (n_1464));
XOR2_X1 i_97 (.Z (n_4729), .A (n_4727), .B (n_436));
AOI21_X1 i_96 (.ZN (n_435), .A (n_4728), .B1 (n_4727), .B2 (n_436));
INV_X1 i_95 (.ZN (n_4731), .A (n_435));
XNOR2_X1 i_94 (.ZN (n_434), .A (n_4855), .B (n_1336));
XOR2_X1 i_93 (.Z (n_4862), .A (n_4860), .B (n_434));
AOI21_X1 i_92 (.ZN (n_433), .A (n_4861), .B1 (n_4860), .B2 (n_434));
INV_X1 i_91 (.ZN (n_4864), .A (n_433));
XNOR2_X1 i_90 (.ZN (n_432), .A (n_4983), .B (n_1218));
XOR2_X1 i_89 (.Z (n_4990), .A (n_4988), .B (n_432));
AOI21_X1 i_88 (.ZN (n_431), .A (n_4989), .B1 (n_4988), .B2 (n_432));
INV_X1 i_87 (.ZN (n_4992), .A (n_431));
XOR2_X1 i_86 (.Z (n_430), .A (n_5103), .B (n_1109));
XOR2_X1 i_85 (.Z (n_5110), .A (n_5108), .B (n_430));
AOI21_X1 i_84 (.ZN (n_429), .A (n_5109), .B1 (n_5108), .B2 (n_430));
INV_X1 i_83 (.ZN (n_5112), .A (n_429));
XNOR2_X1 i_82 (.ZN (n_428), .A (n_5219), .B (n_1014));
XOR2_X1 i_81 (.Z (n_5226), .A (n_5224), .B (n_428));
AOI21_X1 i_80 (.ZN (n_427), .A (n_5225), .B1 (n_5224), .B2 (n_428));
INV_X1 i_79 (.ZN (n_5228), .A (n_427));
XNOR2_X1 i_78 (.ZN (n_426), .A (n_5330), .B (n_954));
XOR2_X1 i_77 (.Z (n_5337), .A (n_5335), .B (n_426));
AOI21_X1 i_76 (.ZN (n_425), .A (n_5336), .B1 (n_5335), .B2 (n_426));
INV_X1 i_75 (.ZN (n_5339), .A (n_425));
XNOR2_X1 i_74 (.ZN (n_424), .A (n_5433), .B (n_897));
XOR2_X1 i_73 (.Z (n_5440), .A (n_5438), .B (n_424));
AOI21_X1 i_72 (.ZN (n_423), .A (n_5439), .B1 (n_5438), .B2 (n_424));
INV_X1 i_71 (.ZN (n_5442), .A (n_423));
XNOR2_X1 i_70 (.ZN (n_422), .A (n_5532), .B (n_840));
XOR2_X1 i_69 (.Z (n_5539), .A (n_5537), .B (n_422));
AOI21_X1 i_68 (.ZN (n_421), .A (n_5538), .B1 (n_5537), .B2 (n_422));
INV_X1 i_67 (.ZN (n_5541), .A (n_421));
XNOR2_X1 i_66 (.ZN (n_420), .A (n_5626), .B (n_793));
XOR2_X1 i_65 (.Z (n_5633), .A (n_5631), .B (n_420));
AOI21_X1 i_64 (.ZN (n_419), .A (n_5632), .B1 (n_5631), .B2 (n_420));
INV_X1 i_63 (.ZN (n_5635), .A (n_419));
XNOR2_X1 i_62 (.ZN (n_418), .A (n_5712), .B (n_748));
XOR2_X1 i_61 (.Z (n_5719), .A (n_5717), .B (n_418));
AOI21_X1 i_60 (.ZN (n_417), .A (n_5718), .B1 (n_5717), .B2 (n_418));
INV_X1 i_59 (.ZN (n_5721), .A (n_417));
XNOR2_X1 i_58 (.ZN (n_416), .A (n_10), .B (n_700));
XOR2_X1 i_57 (.Z (n_272), .A (n_12), .B (n_416));
XNOR2_X1 i_56 (.ZN (n_415), .A (n_26), .B (n_671));
XOR2_X1 i_55 (.Z (n_271), .A (n_28), .B (n_415));
AOI21_X1 i_54 (.ZN (n_414), .A (n_13), .B1 (n_12), .B2 (n_416));
INV_X1 i_53 (.ZN (n_270), .A (n_414));
AOI21_X1 i_52 (.ZN (n_413), .A (n_29), .B1 (n_28), .B2 (n_415));
INV_X1 i_51 (.ZN (n_269), .A (n_413));
XNOR2_X1 i_50 (.ZN (n_412), .A (n_42), .B (n_624));
XOR2_X1 i_49 (.Z (n_268), .A (n_44), .B (n_412));
AOI21_X1 i_48 (.ZN (n_411), .A (n_45), .B1 (n_44), .B2 (n_412));
INV_X1 i_47 (.ZN (n_267), .A (n_411));
XNOR2_X1 i_46 (.ZN (n_410), .A (n_56), .B (n_590));
XOR2_X1 i_45 (.Z (n_266), .A (n_58), .B (n_410));
XNOR2_X1 i_44 (.ZN (n_409), .A (n_68), .B (n_561));
XOR2_X1 i_43 (.Z (n_265), .A (n_70), .B (n_409));
AOI21_X1 i_42 (.ZN (n_408), .A (n_59), .B1 (n_58), .B2 (n_410));
INV_X1 i_41 (.ZN (n_264), .A (n_408));
AOI21_X1 i_40 (.ZN (n_407), .A (n_71), .B1 (n_70), .B2 (n_409));
INV_X1 i_39 (.ZN (n_263), .A (n_407));
XNOR2_X1 i_38 (.ZN (n_406), .A (n_80), .B (n_535));
XOR2_X1 i_37 (.Z (n_262), .A (n_82), .B (n_406));
AOI21_X1 i_36 (.ZN (n_405), .A (n_83), .B1 (n_82), .B2 (n_406));
INV_X1 i_35 (.ZN (n_261), .A (n_405));
XOR2_X1 i_34 (.Z (n_404), .A (n_88), .B (n_508));
XOR2_X1 i_33 (.Z (n_403), .A (n_90), .B (n_404));
XOR2_X1 i_32 (.Z (n_260), .A (n_92), .B (n_403));
AOI21_X1 i_31 (.ZN (n_402), .A (n_91), .B1 (n_90), .B2 (n_404));
INV_X1 i_30 (.ZN (n_401), .A (n_402));
XNOR2_X1 i_29 (.ZN (n_259), .A (n_100), .B (n_402));
AOI21_X1 i_28 (.ZN (n_400), .A (n_93), .B1 (n_92), .B2 (n_403));
INV_X1 i_27 (.ZN (n_258), .A (n_400));
AOI21_X1 i_26 (.ZN (n_399), .A (n_101), .B1 (n_100), .B2 (n_401));
INV_X1 i_25 (.ZN (n_257), .A (n_399));
XNOR2_X1 i_24 (.ZN (n_398), .A (n_106), .B (n_476));
XOR2_X1 i_23 (.Z (n_256), .A (n_108), .B (n_398));
XOR2_X1 i_22 (.Z (n_397), .A (n_112), .B (n_465));
XOR2_X1 i_21 (.Z (n_255), .A (n_114), .B (n_397));
AOI21_X1 i_20 (.ZN (n_396), .A (n_109), .B1 (n_108), .B2 (n_398));
INV_X1 i_19 (.ZN (n_254), .A (n_396));
AOI21_X1 i_18 (.ZN (n_395), .A (n_115), .B1 (n_114), .B2 (n_397));
INV_X1 i_17 (.ZN (n_253), .A (n_395));
OAI21_X1 i_16 (.ZN (n_394), .A (n_461), .B1 (n_484), .B2 (n_462));
XOR2_X1 i_15 (.Z (n_393), .A (n_460), .B (n_394));
XOR2_X1 i_14 (.Z (n_392), .A (n_116), .B (n_393));
XOR2_X1 i_13 (.Z (n_252), .A (n_118), .B (n_392));
AOI21_X1 i_12 (.ZN (n_391), .A (n_117), .B1 (n_116), .B2 (n_393));
INV_X1 i_11 (.ZN (n_390), .A (n_391));
XNOR2_X1 i_10 (.ZN (n_251), .A (n_122), .B (n_391));
AOI21_X1 i_9 (.ZN (n_389), .A (n_119), .B1 (n_118), .B2 (n_392));
INV_X1 i_8 (.ZN (n_250), .A (n_389));
AOI21_X1 i_7 (.ZN (n_388), .A (n_123), .B1 (n_122), .B2 (n_390));
INV_X1 i_6 (.ZN (n_249), .A (n_388));
AOI21_X1 i_5 (.ZN (n_387), .A (n_121), .B1 (n_120), .B2 (n_454));
INV_X1 i_4 (.ZN (n_386), .A (n_387));
XNOR2_X1 i_3 (.ZN (n_248), .A (n_124), .B (n_387));
XOR2_X1 i_2 (.Z (n_247), .A (n_126), .B (n_5742));
AOI21_X1 i_1 (.ZN (n_385), .A (n_125), .B1 (n_124), .B2 (n_386));
INV_X1 i_0 (.ZN (n_246), .A (n_385));
HA_X1 i_6010 (.CO (n_245), .S (n_244), .A (n_247), .B (n_246));
HA_X1 i_6006 (.CO (n_243), .S (n_242), .A (n_249), .B (n_248));
HA_X1 i_6002 (.CO (n_241), .S (n_240), .A (n_251), .B (n_250));
HA_X1 i_5998 (.CO (n_239), .S (n_238), .A (n_253), .B (n_252));
HA_X1 i_5994 (.CO (n_237), .S (n_236), .A (n_255), .B (n_254));
HA_X1 i_5990 (.CO (n_235), .S (n_234), .A (n_257), .B (n_256));
HA_X1 i_5986 (.CO (n_233), .S (n_232), .A (n_259), .B (n_258));
HA_X1 i_5982 (.CO (n_231), .S (n_230), .A (n_261), .B (n_260));
HA_X1 i_5978 (.CO (n_229), .S (n_228), .A (n_263), .B (n_262));
HA_X1 i_5974 (.CO (n_227), .S (n_226), .A (n_265), .B (n_264));
HA_X1 i_5970 (.CO (n_225), .S (n_224), .A (n_267), .B (n_266));
HA_X1 i_5966 (.CO (n_223), .S (n_222), .A (n_269), .B (n_268));
HA_X1 i_5962 (.CO (n_221), .S (n_220), .A (n_271), .B (n_270));
HA_X1 i_5958 (.CO (n_219), .S (n_218), .A (n_5721), .B (n_272));
HA_X1 i_5954 (.CO (n_217), .S (n_216), .A (n_5635), .B (n_5719));
HA_X1 i_5950 (.CO (n_215), .S (n_214), .A (n_5541), .B (n_5633));
HA_X1 i_5946 (.CO (n_213), .S (n_212), .A (n_5442), .B (n_5539));
HA_X1 i_5942 (.CO (n_211), .S (n_210), .A (n_5339), .B (n_5440));
HA_X1 i_5938 (.CO (n_209), .S (n_208), .A (n_5228), .B (n_5337));
HA_X1 i_5934 (.CO (n_207), .S (n_206), .A (n_5112), .B (n_5226));
HA_X1 i_5930 (.CO (n_205), .S (n_204), .A (n_4992), .B (n_5110));
HA_X1 i_5926 (.CO (n_203), .S (n_202), .A (n_4864), .B (n_4990));
HA_X1 i_5922 (.CO (n_201), .S (n_200), .A (n_4731), .B (n_4862));
HA_X1 i_5918 (.CO (n_199), .S (n_198), .A (n_4594), .B (n_4729));
HA_X1 i_5914 (.CO (n_197), .S (n_196), .A (n_4449), .B (n_4592));
HA_X1 i_5910 (.CO (n_195), .S (n_194), .A (n_4299), .B (n_4447));
HA_X1 i_5906 (.CO (n_193), .S (n_192), .A (n_4297), .B (n_4145));
HA_X1 i_5902 (.CO (n_191), .S (n_190), .A (n_3983), .B (n_4143));
HA_X1 i_5898 (.CO (n_189), .S (n_188), .A (n_3816), .B (n_3981));
HA_X1 i_5894 (.CO (n_187), .S (n_186), .A (n_3646), .B (n_3814));
HA_X1 i_5890 (.CO (n_185), .S (n_184), .A (n_3475), .B (n_3645));
HA_X1 i_5886 (.CO (n_183), .S (n_182), .A (n_3310), .B (n_3474));
HA_X1 i_5882 (.CO (n_181), .S (n_180), .A (n_3153), .B (n_3309));
HA_X1 i_5878 (.CO (n_179), .S (n_178), .A (n_3000), .B (n_3152));
HA_X1 i_5874 (.CO (n_177), .S (n_176), .A (n_2852), .B (n_2999));
HA_X1 i_5870 (.CO (n_175), .S (n_174), .A (n_2712), .B (n_2851));
HA_X1 i_5866 (.CO (n_173), .S (n_172), .A (n_2708), .B (n_2711));
HA_X1 i_5862 (.CO (n_171), .S (n_170), .A (n_2445), .B (n_2575));
HA_X1 i_5858 (.CO (n_169), .S (n_168), .A (n_2322), .B (n_2444));
HA_X1 i_5854 (.CO (n_167), .S (n_166), .A (n_2203), .B (n_2321));
HA_X1 i_5850 (.CO (n_165), .S (n_164), .A (n_2089), .B (n_2202));
HA_X1 i_5846 (.CO (n_163), .S (n_162), .A (n_2085), .B (n_2088));
HA_X1 i_5842 (.CO (n_161), .S (n_160), .A (n_1881), .B (n_1982));
HA_X1 i_5838 (.CO (n_159), .S (n_158), .A (n_1784), .B (n_1880));
HA_X1 i_5834 (.CO (n_157), .S (n_156), .A (n_1780), .B (n_1783));
HA_X1 i_5830 (.CO (n_155), .S (n_154), .A (n_1691), .B (n_1694));
HA_X1 i_5826 (.CO (n_153), .S (n_152), .A (n_1606), .B (n_1609));
HA_X1 i_5822 (.CO (n_151), .S (n_150), .A (n_1526), .B (n_1529));
HA_X1 i_5818 (.CO (n_149), .S (n_148), .A (n_1454), .B (n_1457));
HA_X1 i_5814 (.CO (n_147), .S (n_146), .A (n_1386), .B (n_1389));
HA_X1 i_5810 (.CO (n_145), .S (n_144), .A (n_1323), .B (n_1326));
HA_X1 i_5806 (.CO (n_143), .S (n_142), .A (n_1271), .B (n_1268));
HA_X1 i_5802 (.CO (n_141), .S (n_140), .A (n_1220), .B (n_1217));
HA_X1 i_5798 (.CO (n_139), .S (n_138), .A (n_1171), .B (n_1174));
HA_X1 i_5794 (.CO (n_137), .S (n_136), .A (n_1133), .B (n_1136));
HA_X1 i_5790 (.CO (n_135), .S (n_134), .A (n_1102), .B (n_1099));
HA_X1 i_5786 (.CO (n_133), .S (n_132), .A (n_1073), .B (n_1070));
HA_X1 i_5782 (.CO (n_131), .S (n_130), .A (n_1039), .B (n_1052));
HA_X1 i_5778 (.CO (n_129), .S (n_128), .A (n_1034), .B (n_1029));
HA_X1 i_5762 (.CO (n_127), .S (n_126), .A (n_1022), .B (n_991));
HA_X1 i_5758 (.CO (n_125), .S (n_124), .A (n_274), .B (n_273));
HA_X1 i_5746 (.CO (n_123), .S (n_122), .A (n_276), .B (n_275));
HA_X1 i_5742 (.CO (n_121), .S (n_120), .A (n_927), .B (n_277));
HA_X1 i_5730 (.CO (n_119), .S (n_118), .A (n_279), .B (n_278));
HA_X1 i_5726 (.CO (n_117), .S (n_116), .A (n_281), .B (n_280));
HA_X1 i_5706 (.CO (n_115), .S (n_114), .A (n_283), .B (n_282));
HA_X1 i_5702 (.CO (n_113), .S (n_112), .A (n_285), .B (n_284));
HA_X1 i_5698 (.CO (n_111), .S (n_110), .A (n_287), .B (n_286));
HA_X1 i_5678 (.CO (n_109), .S (n_108), .A (n_289), .B (n_288));
HA_X1 i_5674 (.CO (n_107), .S (n_106), .A (n_291), .B (n_290));
HA_X1 i_5670 (.CO (n_105), .S (n_104), .A (n_293), .B (n_292));
HA_X1 i_5666 (.CO (n_103), .S (n_102), .A (n_831), .B (n_294));
HA_X1 i_5647 (.CO (n_101), .S (n_100), .A (n_296), .B (n_295));
HA_X1 i_5643 (.CO (n_99), .S (n_98), .A (n_298), .B (n_297));
HA_X1 i_5639 (.CO (n_97), .S (n_96), .A (n_300), .B (n_299));
HA_X1 i_5635 (.CO (n_95), .S (n_94), .A (n_302), .B (n_301));
HA_X1 i_5608 (.CO (n_93), .S (n_92), .A (n_304), .B (n_303));
HA_X1 i_5604 (.CO (n_91), .S (n_90), .A (n_306), .B (n_305));
HA_X1 i_5600 (.CO (n_89), .S (n_88), .A (n_308), .B (n_307));
HA_X1 i_5596 (.CO (n_87), .S (n_86), .A (n_310), .B (n_309));
HA_X1 i_5592 (.CO (n_85), .S (n_84), .A (n_312), .B (n_311));
HA_X1 i_5565 (.CO (n_83), .S (n_82), .A (n_314), .B (n_313));
HA_X1 i_5561 (.CO (n_81), .S (n_80), .A (n_316), .B (n_315));
HA_X1 i_5557 (.CO (n_79), .S (n_78), .A (n_318), .B (n_317));
HA_X1 i_5553 (.CO (n_77), .S (n_76), .A (n_320), .B (n_319));
HA_X1 i_5549 (.CO (n_75), .S (n_74), .A (n_322), .B (n_321));
HA_X1 i_5545 (.CO (n_73), .S (n_72), .A (n_735), .B (n_323));
HA_X1 i_5519 (.CO (n_71), .S (n_70), .A (n_325), .B (n_324));
HA_X1 i_5515 (.CO (n_69), .S (n_68), .A (n_327), .B (n_326));
HA_X1 i_5511 (.CO (n_67), .S (n_66), .A (n_329), .B (n_328));
HA_X1 i_5507 (.CO (n_65), .S (n_64), .A (n_331), .B (n_330));
HA_X1 i_5503 (.CO (n_63), .S (n_62), .A (n_333), .B (n_332));
HA_X1 i_5499 (.CO (n_61), .S (n_60), .A (n_335), .B (n_334));
HA_X1 i_5465 (.CO (n_59), .S (n_58), .A (n_337), .B (n_336));
HA_X1 i_5461 (.CO (n_57), .S (n_56), .A (n_339), .B (n_338));
HA_X1 i_5457 (.CO (n_55), .S (n_54), .A (n_341), .B (n_340));
HA_X1 i_5453 (.CO (n_53), .S (n_52), .A (n_343), .B (n_342));
HA_X1 i_5449 (.CO (n_51), .S (n_50), .A (n_345), .B (n_344));
HA_X1 i_5445 (.CO (n_49), .S (n_48), .A (n_347), .B (n_346));
HA_X1 i_5441 (.CO (n_47), .S (n_46), .A (n_349), .B (n_348));
HA_X1 i_5407 (.CO (n_45), .S (n_44), .A (n_351), .B (n_350));
HA_X1 i_5403 (.CO (n_43), .S (n_42), .A (n_353), .B (n_352));
HA_X1 i_5399 (.CO (n_41), .S (n_40), .A (n_355), .B (n_354));
HA_X1 i_5395 (.CO (n_39), .S (n_38), .A (n_357), .B (n_356));
HA_X1 i_5391 (.CO (n_37), .S (n_36), .A (n_359), .B (n_358));
HA_X1 i_5387 (.CO (n_35), .S (n_34), .A (n_361), .B (n_360));
HA_X1 i_5383 (.CO (n_33), .S (n_32), .A (n_363), .B (n_362));
HA_X1 i_5379 (.CO (n_31), .S (n_30), .A (n_639), .B (n_364));
HA_X1 i_5346 (.CO (n_29), .S (n_28), .A (n_366), .B (n_365));
HA_X1 i_5342 (.CO (n_27), .S (n_26), .A (n_368), .B (n_367));
HA_X1 i_5338 (.CO (n_25), .S (n_24), .A (n_370), .B (n_369));
HA_X1 i_5334 (.CO (n_23), .S (n_22), .A (n_372), .B (n_371));
HA_X1 i_5330 (.CO (n_21), .S (n_20), .A (n_374), .B (n_373));
HA_X1 i_5326 (.CO (n_19), .S (n_18), .A (n_376), .B (n_375));
HA_X1 i_5322 (.CO (n_17), .S (n_16), .A (n_5724), .B (n_5763));
HA_X1 i_5318 (.CO (n_15), .S (n_14), .A (n_5747), .B (n_5740));
HA_X1 i_5277 (.CO (n_13), .S (n_12), .A (n_377), .B (n_5716));
HA_X1 i_5273 (.CO (n_11), .S (n_10), .A (n_379), .B (n_378));
HA_X1 i_5269 (.CO (n_9), .S (n_8), .A (n_381), .B (n_380));
HA_X1 i_5265 (.CO (n_7), .S (n_6), .A (n_5686), .B (n_5701));
HA_X1 i_5261 (.CO (n_5), .S (n_4), .A (n_5766), .B (n_5761));
HA_X1 i_5257 (.CO (n_3), .S (n_2), .A (n_5739), .B (n_5732));
HA_X1 i_5253 (.CO (n_1), .S (n_0), .A (n_5676), .B (n_5752));
HA_X1 i_5249 (.CO (n_5765), .S (n_5764), .A (n_5647), .B (n_5638));
HA_X1 i_5245 (.CO (n_5760), .S (n_5759), .A (n_5668), .B (n_5661));
HA_X1 i_5204 (.CO (n_5718), .S (n_5717), .A (n_5709), .B (n_5630));
HA_X1 i_5200 (.CO (n_5713), .S (n_5712), .A (n_5620), .B (n_5704));
HA_X1 i_5196 (.CO (n_5708), .S (n_5707), .A (n_5689), .B (n_5694));
HA_X1 i_5192 (.CO (n_5703), .S (n_5702), .A (n_5684), .B (n_5610));
HA_X1 i_5188 (.CO (n_5698), .S (n_5697), .A (n_5674), .B (n_5605));
HA_X1 i_5184 (.CO (n_5693), .S (n_5692), .A (n_5637), .B (n_5595));
HA_X1 i_5180 (.CO (n_5688), .S (n_5687), .A (n_5660), .B (n_5653));
HA_X1 i_5176 (.CO (n_5683), .S (n_5682), .A (n_5590), .B (n_5581));
HA_X1 i_5172 (.CO (n_5678), .S (n_5677), .A (n_5560), .B (n_5553));
HA_X1 i_5168 (.CO (n_5673), .S (n_5672), .A (n_543), .B (n_5574));
HA_X1 i_5128 (.CO (n_5632), .S (n_5631), .A (n_5623), .B (n_5536));
HA_X1 i_5124 (.CO (n_5627), .S (n_5626), .A (n_5526), .B (n_5618));
HA_X1 i_5120 (.CO (n_5622), .S (n_5621), .A (n_5521), .B (n_5613));
HA_X1 i_5116 (.CO (n_5617), .S (n_5616), .A (n_5516), .B (n_5603));
HA_X1 i_5112 (.CO (n_5612), .S (n_5611), .A (n_5506), .B (n_5501));
HA_X1 i_5108 (.CO (n_5607), .S (n_5606), .A (n_5543), .B (n_5593));
HA_X1 i_5104 (.CO (n_5602), .S (n_5601), .A (n_5566), .B (n_5559));
HA_X1 i_5100 (.CO (n_5597), .S (n_5596), .A (n_5491), .B (n_5580));
HA_X1 i_5096 (.CO (n_5592), .S (n_5591), .A (n_5454), .B (n_5445));
HA_X1 i_5092 (.CO (n_5587), .S (n_5586), .A (n_5475), .B (n_5468));
HA_X1 i_5044 (.CO (n_5538), .S (n_5537), .A (n_5529), .B (n_5437));
HA_X1 i_5040 (.CO (n_5533), .S (n_5532), .A (n_5427), .B (n_5524));
HA_X1 i_5036 (.CO (n_5528), .S (n_5527), .A (n_5514), .B (n_5422));
HA_X1 i_5032 (.CO (n_5523), .S (n_5522), .A (n_5412), .B (n_5509));
HA_X1 i_5028 (.CO (n_5518), .S (n_5517), .A (n_5402), .B (n_5499));
HA_X1 i_5024 (.CO (n_5513), .S (n_5512), .A (n_5494), .B (n_5489));
HA_X1 i_5020 (.CO (n_5508), .S (n_5507), .A (n_5453), .B (n_5444));
HA_X1 i_5016 (.CO (n_5503), .S (n_5502), .A (n_5474), .B (n_5467));
HA_X1 i_5012 (.CO (n_5498), .S (n_5497), .A (n_5392), .B (n_5387));
HA_X1 i_5008 (.CO (n_5493), .S (n_5492), .A (n_5358), .B (n_5351));
HA_X1 i_5004 (.CO (n_5488), .S (n_5487), .A (n_5379), .B (n_5372));
HA_X1 i_4956 (.CO (n_5439), .S (n_5438), .A (n_5430), .B (n_5334));
HA_X1 i_4952 (.CO (n_5434), .S (n_5433), .A (n_5324), .B (n_5425));
HA_X1 i_4948 (.CO (n_5429), .S (n_5428), .A (n_5410), .B (n_5319));
HA_X1 i_4944 (.CO (n_5424), .S (n_5423), .A (n_5400), .B (n_5314));
HA_X1 i_4940 (.CO (n_5419), .S (n_5418), .A (n_5395), .B (n_5309));
HA_X1 i_4936 (.CO (n_5414), .S (n_5413), .A (n_5304), .B (n_5299));
HA_X1 i_4932 (.CO (n_5409), .S (n_5408), .A (n_5341), .B (n_5390));
HA_X1 i_4928 (.CO (n_5404), .S (n_5403), .A (n_5364), .B (n_5357));
HA_X1 i_4924 (.CO (n_5399), .S (n_5398), .A (n_5275), .B (n_5378));
HA_X1 i_4920 (.CO (n_5394), .S (n_5393), .A (n_5231), .B (n_5289));
HA_X1 i_4916 (.CO (n_5389), .S (n_5388), .A (n_5254), .B (n_5247));
HA_X1 i_4912 (.CO (n_5384), .S (n_5383), .A (n_447), .B (n_5268));
HA_X1 i_4865 (.CO (n_5336), .S (n_5335), .A (n_5327), .B (n_5223));
HA_X1 i_4861 (.CO (n_5331), .S (n_5330), .A (n_5213), .B (n_5322));
HA_X1 i_4857 (.CO (n_5326), .S (n_5325), .A (n_5307), .B (n_5208));
HA_X1 i_4853 (.CO (n_5321), .S (n_5320), .A (n_5297), .B (n_5203));
HA_X1 i_4849 (.CO (n_5316), .S (n_5315), .A (n_5198), .B (n_5193));
HA_X1 i_4845 (.CO (n_5311), .S (n_5310), .A (n_5188), .B (n_5183));
HA_X1 i_4841 (.CO (n_5306), .S (n_5305), .A (n_5178), .B (n_5287));
HA_X1 i_4837 (.CO (n_5301), .S (n_5300), .A (n_5246), .B (n_5239));
HA_X1 i_4833 (.CO (n_5296), .S (n_5295), .A (n_5267), .B (n_5260));
HA_X1 i_4829 (.CO (n_5291), .S (n_5290), .A (n_5173), .B (n_5168));
HA_X1 i_4825 (.CO (n_5286), .S (n_5285), .A (n_5131), .B (n_5124));
HA_X1 i_4821 (.CO (n_5281), .S (n_5280), .A (n_5152), .B (n_5145));
HA_X1 i_4766 (.CO (n_5225), .S (n_5224), .A (n_5216), .B (n_5107));
HA_X1 i_4762 (.CO (n_5220), .S (n_5219), .A (n_5206), .B (n_5211));
HA_X1 i_4758 (.CO (n_5215), .S (n_5214), .A (n_5092), .B (n_5201));
HA_X1 i_4754 (.CO (n_5210), .S (n_5209), .A (n_5191), .B (n_5087));
HA_X1 i_4750 (.CO (n_5205), .S (n_5204), .A (n_5077), .B (n_5186));
HA_X1 i_4746 (.CO (n_5200), .S (n_5199), .A (n_5062), .B (n_5176));
HA_X1 i_4742 (.CO (n_5195), .S (n_5194), .A (n_5166), .B (n_5072));
HA_X1 i_4738 (.CO (n_5190), .S (n_5189), .A (n_5114), .B (n_5057));
HA_X1 i_4734 (.CO (n_5185), .S (n_5184), .A (n_5137), .B (n_5130));
HA_X1 i_4730 (.CO (n_5180), .S (n_5179), .A (n_5157), .B (n_5151));
HA_X1 i_4726 (.CO (n_5175), .S (n_5174), .A (n_4995), .B (n_5052));
HA_X1 i_4722 (.CO (n_5170), .S (n_5169), .A (n_5018), .B (n_5011));
HA_X1 i_4718 (.CO (n_5165), .S (n_5164), .A (n_5039), .B (n_5032));
HA_X1 i_4663 (.CO (n_5109), .S (n_5108), .A (n_5100), .B (n_4987));
HA_X1 i_4659 (.CO (n_5104), .S (n_5103), .A (n_5090), .B (n_4982));
HA_X1 i_4655 (.CO (n_5099), .S (n_5098), .A (n_4972), .B (n_5085));
HA_X1 i_4651 (.CO (n_5094), .S (n_5093), .A (n_5080), .B (n_5075));
HA_X1 i_4647 (.CO (n_5089), .S (n_5088), .A (n_5070), .B (n_5065));
HA_X1 i_4643 (.CO (n_5084), .S (n_5083), .A (n_4952), .B (n_5060));
HA_X1 i_4639 (.CO (n_5079), .S (n_5078), .A (n_5045), .B (n_4947));
HA_X1 i_4635 (.CO (n_5074), .S (n_5073), .A (n_4937), .B (n_5055));
HA_X1 i_4631 (.CO (n_5069), .S (n_5068), .A (n_5010), .B (n_5003));
HA_X1 i_4627 (.CO (n_5064), .S (n_5063), .A (n_5031), .B (n_5024));
HA_X1 i_4623 (.CO (n_5059), .S (n_5058), .A (n_4927), .B (n_4918));
HA_X1 i_4619 (.CO (n_5054), .S (n_5053), .A (n_4876), .B (n_4867));
HA_X1 i_4615 (.CO (n_5049), .S (n_5048), .A (n_4897), .B (n_4890));
HA_X1 i_4611 (.CO (n_5044), .S (n_5043), .A (n_382), .B (n_4911));
HA_X1 i_4557 (.CO (n_4989), .S (n_4988), .A (n_4980), .B (n_4859));
HA_X1 i_4553 (.CO (n_4984), .S (n_4983), .A (n_4970), .B (n_4975));
HA_X1 i_4549 (.CO (n_4979), .S (n_4978), .A (n_4844), .B (n_4965));
HA_X1 i_4545 (.CO (n_4974), .S (n_4973), .A (n_4960), .B (n_4955));
HA_X1 i_4541 (.CO (n_4969), .S (n_4968), .A (n_4945), .B (n_4940));
HA_X1 i_4537 (.CO (n_4964), .S (n_4963), .A (n_4829), .B (n_4824));
HA_X1 i_4533 (.CO (n_4959), .S (n_4958), .A (n_4814), .B (n_4809));
HA_X1 i_4529 (.CO (n_4954), .S (n_4953), .A (n_4930), .B (n_4925));
HA_X1 i_4525 (.CO (n_4949), .S (n_4948), .A (n_4875), .B (n_4866));
HA_X1 i_4521 (.CO (n_4944), .S (n_4943), .A (n_4896), .B (n_4889));
HA_X1 i_4517 (.CO (n_4939), .S (n_4938), .A (n_4917), .B (n_4910));
HA_X1 i_4513 (.CO (n_4934), .S (n_4933), .A (n_4734), .B (n_4799));
HA_X1 i_4509 (.CO (n_4929), .S (n_4928), .A (n_4757), .B (n_4750));
HA_X1 i_4505 (.CO (n_4924), .S (n_4923), .A (n_4778), .B (n_4771));
HA_X1 i_4443 (.CO (n_4861), .S (n_4860), .A (n_4852), .B (n_4726));
HA_X1 i_4439 (.CO (n_4856), .S (n_4855), .A (n_4716), .B (n_4847));
HA_X1 i_4435 (.CO (n_4851), .S (n_4850), .A (n_4837), .B (n_4711));
HA_X1 i_4431 (.CO (n_4846), .S (n_4845), .A (n_4827), .B (n_4706));
HA_X1 i_4427 (.CO (n_4841), .S (n_4840), .A (n_4812), .B (n_4822));
HA_X1 i_4423 (.CO (n_4836), .S (n_4835), .A (n_4696), .B (n_4691));
HA_X1 i_4419 (.CO (n_4831), .S (n_4830), .A (n_4676), .B (n_4686));
HA_X1 i_4415 (.CO (n_4826), .S (n_4825), .A (n_4797), .B (n_4792));
HA_X1 i_4411 (.CO (n_4821), .S (n_4820), .A (n_4733), .B (n_4671));
HA_X1 i_4407 (.CO (n_4816), .S (n_4815), .A (n_4756), .B (n_4749));
HA_X1 i_4403 (.CO (n_4811), .S (n_4810), .A (n_4777), .B (n_4770));
HA_X1 i_4399 (.CO (n_4806), .S (n_4805), .A (n_4661), .B (n_4656));
HA_X1 i_4395 (.CO (n_4801), .S (n_4800), .A (n_4606), .B (n_4597));
HA_X1 i_4391 (.CO (n_4796), .S (n_4795), .A (n_4627), .B (n_4620));
HA_X1 i_4387 (.CO (n_4791), .S (n_4790), .A (n_4648), .B (n_4641));
HA_X1 i_4325 (.CO (n_4728), .S (n_4727), .A (n_4589), .B (n_4719));
HA_X1 i_4321 (.CO (n_4723), .S (n_4722), .A (n_4579), .B (n_4714));
HA_X1 i_4317 (.CO (n_4718), .S (n_4717), .A (n_4574), .B (n_4704));
HA_X1 i_4313 (.CO (n_4713), .S (n_4712), .A (n_4689), .B (n_4569));
HA_X1 i_4309 (.CO (n_4708), .S (n_4707), .A (n_4674), .B (n_4564));
HA_X1 i_4305 (.CO (n_4703), .S (n_4702), .A (n_4554), .B (n_4684));
HA_X1 i_4301 (.CO (n_4698), .S (n_4697), .A (n_4549), .B (n_4669));
HA_X1 i_4297 (.CO (n_4693), .S (n_4692), .A (n_4544), .B (n_4539));
HA_X1 i_4293 (.CO (n_4688), .S (n_4687), .A (n_4664), .B (n_4659));
HA_X1 i_4289 (.CO (n_4683), .S (n_4682), .A (n_4605), .B (n_4596));
HA_X1 i_4285 (.CO (n_4678), .S (n_4677), .A (n_4626), .B (n_4619));
HA_X1 i_4281 (.CO (n_4673), .S (n_4672), .A (n_4647), .B (n_4640));
HA_X1 i_4277 (.CO (n_4668), .S (n_4667), .A (n_4524), .B (n_4519));
HA_X1 i_4273 (.CO (n_4663), .S (n_4662), .A (n_4468), .B (n_4461));
HA_X1 i_4269 (.CO (n_4658), .S (n_4657), .A (n_4489), .B (n_4482));
HA_X1 i_4265 (.CO (n_4653), .S (n_4652), .A (n_383), .B (n_4503));
HA_X1 i_4204 (.CO (n_4591), .S (n_4590), .A (n_4444), .B (n_4582));
HA_X1 i_4200 (.CO (n_4586), .S (n_4585), .A (n_4572), .B (n_4577));
HA_X1 i_4196 (.CO (n_4581), .S (n_4580), .A (n_4429), .B (n_4567));
HA_X1 i_4192 (.CO (n_4576), .S (n_4575), .A (n_4419), .B (n_4424));
HA_X1 i_4188 (.CO (n_4571), .S (n_4570), .A (n_4414), .B (n_4557));
HA_X1 i_4184 (.CO (n_4566), .S (n_4565), .A (n_4547), .B (n_4542));
HA_X1 i_4180 (.CO (n_4561), .S (n_4560), .A (n_4532), .B (n_4409));
HA_X1 i_4176 (.CO (n_4556), .S (n_4555), .A (n_4399), .B (n_4394));
HA_X1 i_4172 (.CO (n_4551), .S (n_4550), .A (n_4527), .B (n_4522));
HA_X1 i_4168 (.CO (n_4546), .S (n_4545), .A (n_4460), .B (n_4451));
HA_X1 i_4164 (.CO (n_4541), .S (n_4540), .A (n_4481), .B (n_4474));
HA_X1 i_4160 (.CO (n_4536), .S (n_4535), .A (n_4502), .B (n_4495));
HA_X1 i_4156 (.CO (n_4531), .S (n_4530), .A (n_4374), .B (n_4369));
HA_X1 i_4152 (.CO (n_4526), .S (n_4525), .A (n_4311), .B (n_4302));
HA_X1 i_4148 (.CO (n_4521), .S (n_4520), .A (n_4332), .B (n_4325));
HA_X1 i_4144 (.CO (n_4516), .S (n_4515), .A (n_4353), .B (n_4346));
HA_X1 i_4075 (.CO (n_4446), .S (n_4445), .A (n_4437), .B (n_4294));
HA_X1 i_4071 (.CO (n_4441), .S (n_4440), .A (n_4427), .B (n_4432));
HA_X1 i_4067 (.CO (n_4436), .S (n_4435), .A (n_4279), .B (n_4422));
HA_X1 i_4063 (.CO (n_4431), .S (n_4430), .A (n_4412), .B (n_4274));
HA_X1 i_4059 (.CO (n_4426), .S (n_4425), .A (n_4407), .B (n_4402));
HA_X1 i_4055 (.CO (n_4421), .S (n_4420), .A (n_4392), .B (n_4387));
HA_X1 i_4051 (.CO (n_4416), .S (n_4415), .A (n_4259), .B (n_4254));
HA_X1 i_4047 (.CO (n_4411), .S (n_4410), .A (n_4234), .B (n_4249));
HA_X1 i_4043 (.CO (n_4406), .S (n_4405), .A (n_4367), .B (n_4244));
HA_X1 i_4039 (.CO (n_4401), .S (n_4400), .A (n_4229), .B (n_4377));
HA_X1 i_4035 (.CO (n_4396), .S (n_4395), .A (n_4317), .B (n_4310));
HA_X1 i_4031 (.CO (n_4391), .S (n_4390), .A (n_4338), .B (n_4331));
HA_X1 i_4027 (.CO (n_4386), .S (n_4385), .A (n_4358), .B (n_4352));
HA_X1 i_4023 (.CO (n_4381), .S (n_4380), .A (n_4224), .B (n_4219));
HA_X1 i_4019 (.CO (n_4376), .S (n_4375), .A (n_4164), .B (n_4157));
HA_X1 i_4015 (.CO (n_4371), .S (n_4370), .A (n_4185), .B (n_4178));
HA_X1 i_4011 (.CO (n_4366), .S (n_4365), .A (n_4206), .B (n_4199));
HA_X1 i_3942 (.CO (n_4296), .S (n_4295), .A (n_4287), .B (n_4140));
HA_X1 i_3938 (.CO (n_4291), .S (n_4290), .A (n_4277), .B (n_4135));
HA_X1 i_3934 (.CO (n_4286), .S (n_4285), .A (n_4125), .B (n_4272));
HA_X1 i_3930 (.CO (n_4281), .S (n_4280), .A (n_4120), .B (n_4267));
HA_X1 i_3926 (.CO (n_4276), .S (n_4275), .A (n_4257), .B (n_4252));
HA_X1 i_3922 (.CO (n_4271), .S (n_4270), .A (n_4242), .B (n_4237));
HA_X1 i_3918 (.CO (n_4266), .S (n_4265), .A (n_4100), .B (n_4095));
HA_X1 i_3914 (.CO (n_4261), .S (n_4260), .A (n_4232), .B (n_4227));
HA_X1 i_3910 (.CO (n_4256), .S (n_4255), .A (n_4090), .B (n_4085));
HA_X1 i_3906 (.CO (n_4251), .S (n_4250), .A (n_4222), .B (n_4217));
HA_X1 i_3902 (.CO (n_4246), .S (n_4245), .A (n_4156), .B (n_4147));
HA_X1 i_3898 (.CO (n_4241), .S (n_4240), .A (n_4177), .B (n_4170));
HA_X1 i_3894 (.CO (n_4236), .S (n_4235), .A (n_4198), .B (n_4191));
HA_X1 i_3890 (.CO (n_4231), .S (n_4230), .A (n_4060), .B (n_4051));
HA_X1 i_3886 (.CO (n_4226), .S (n_4225), .A (n_3986), .B (n_4070));
HA_X1 i_3882 (.CO (n_4221), .S (n_4220), .A (n_4009), .B (n_4002));
HA_X1 i_3878 (.CO (n_4216), .S (n_4215), .A (n_4030), .B (n_4023));
HA_X1 i_3874 (.CO (n_4211), .S (n_4210), .A (n_384), .B (n_4044));
HA_X1 i_3806 (.CO (n_4142), .S (n_4141), .A (n_4133), .B (n_3978));
HA_X1 i_3802 (.CO (n_4137), .S (n_4136), .A (n_4123), .B (n_4128));
HA_X1 i_3798 (.CO (n_4132), .S (n_4131), .A (n_4113), .B (n_4118));
HA_X1 i_3794 (.CO (n_4127), .S (n_4126), .A (n_4108), .B (n_3963));
HA_X1 i_3790 (.CO (n_4122), .S (n_4121), .A (n_4103), .B (n_4098));
HA_X1 i_3786 (.CO (n_4117), .S (n_4116), .A (n_4093), .B (n_3948));
HA_X1 i_3782 (.CO (n_4112), .S (n_4111), .A (n_4088), .B (n_4083));
HA_X1 i_3778 (.CO (n_4107), .S (n_4106), .A (n_4073), .B (n_3938));
HA_X1 i_3774 (.CO (n_4102), .S (n_4101), .A (n_3923), .B (n_3918));
HA_X1 i_3770 (.CO (n_4097), .S (n_4096), .A (n_4063), .B (n_4058));
HA_X1 i_3766 (.CO (n_4092), .S (n_4091), .A (n_3985), .B (n_3908));
HA_X1 i_3762 (.CO (n_4087), .S (n_4086), .A (n_4008), .B (n_4001));
HA_X1 i_3758 (.CO (n_4082), .S (n_4081), .A (n_4029), .B (n_4022));
HA_X1 i_3754 (.CO (n_4077), .S (n_4076), .A (n_4050), .B (n_4043));
HA_X1 i_3750 (.CO (n_4072), .S (n_4071), .A (n_3903), .B (n_3898));
HA_X1 i_3746 (.CO (n_4067), .S (n_4066), .A (n_3835), .B (n_3828));
HA_X1 i_3742 (.CO (n_4062), .S (n_4061), .A (n_3856), .B (n_3849));
HA_X1 i_3738 (.CO (n_4057), .S (n_4056), .A (n_3877), .B (n_3870));
HA_X1 i_3662 (.CO (n_3980), .S (n_3979), .A (n_3971), .B (n_3811));
HA_X1 i_3658 (.CO (n_3975), .S (n_3974), .A (n_3801), .B (n_3966));
HA_X1 i_3654 (.CO (n_3970), .S (n_3969), .A (n_3951), .B (n_3961));
HA_X1 i_3650 (.CO (n_3965), .S (n_3964), .A (n_3946), .B (n_3791));
HA_X1 i_3646 (.CO (n_3960), .S (n_3959), .A (n_3931), .B (n_3786));
HA_X1 i_3642 (.CO (n_3955), .S (n_3954), .A (n_3776), .B (n_3941));
HA_X1 i_3638 (.CO (n_3950), .S (n_3949), .A (n_3926), .B (n_3921));
HA_X1 i_3634 (.CO (n_3945), .S (n_3944), .A (n_3906), .B (n_3771));
HA_X1 i_3630 (.CO (n_3940), .S (n_3939), .A (n_3751), .B (n_3746));
HA_X1 i_3626 (.CO (n_3935), .S (n_3934), .A (n_3891), .B (n_3761));
HA_X1 i_3622 (.CO (n_3930), .S (n_3929), .A (n_3741), .B (n_3901));
HA_X1 i_3618 (.CO (n_3925), .S (n_3924), .A (n_3834), .B (n_3827));
HA_X1 i_3614 (.CO (n_3920), .S (n_3919), .A (n_3855), .B (n_3848));
HA_X1 i_3610 (.CO (n_3915), .S (n_3914), .A (n_3876), .B (n_3869));
HA_X1 i_3606 (.CO (n_3910), .S (n_3909), .A (n_3726), .B (n_3717));
HA_X1 i_3602 (.CO (n_3905), .S (n_3904), .A (n_3649), .B (n_3736));
HA_X1 i_3598 (.CO (n_3900), .S (n_3899), .A (n_3668), .B (n_3661));
HA_X1 i_3594 (.CO (n_3895), .S (n_3894), .A (n_3689), .B (n_3682));
HA_X1 i_3590 (.CO (n_3890), .S (n_3889), .A (n_3710), .B (n_3703));
HA_X1 i_3514 (.CO (n_3813), .S (n_3812), .A (n_3804), .B (n_3809));
HA_X1 i_3510 (.CO (n_3808), .S (n_3807), .A (n_3634), .B (n_3799));
HA_X1 i_3506 (.CO (n_3803), .S (n_3802), .A (n_3629), .B (n_3789));
HA_X1 i_3502 (.CO (n_3798), .S (n_3797), .A (n_3779), .B (n_3624));
HA_X1 i_3498 (.CO (n_3793), .S (n_3792), .A (n_3614), .B (n_3774));
HA_X1 i_3494 (.CO (n_3788), .S (n_3787), .A (n_3609), .B (n_3769));
HA_X1 i_3490 (.CO (n_3783), .S (n_3782), .A (n_3754), .B (n_3749));
HA_X1 i_3486 (.CO (n_3778), .S (n_3777), .A (n_3604), .B (n_3599));
HA_X1 i_3482 (.CO (n_3773), .S (n_3772), .A (n_3579), .B (n_3594));
HA_X1 i_3478 (.CO (n_3768), .S (n_3767), .A (n_3724), .B (n_3589));
HA_X1 i_3474 (.CO (n_3763), .S (n_3762), .A (n_3574), .B (n_3734));
HA_X1 i_3470 (.CO (n_3758), .S (n_3757), .A (n_3660), .B (n_3653));
HA_X1 i_3466 (.CO (n_3753), .S (n_3752), .A (n_3681), .B (n_3674));
HA_X1 i_3462 (.CO (n_3748), .S (n_3747), .A (n_3702), .B (n_3695));
HA_X1 i_3458 (.CO (n_3743), .S (n_3742), .A (n_3550), .B (n_3716));
HA_X1 i_3454 (.CO (n_3738), .S (n_3737), .A (n_3569), .B (n_3564));
HA_X1 i_3450 (.CO (n_3733), .S (n_3732), .A (n_3494), .B (n_3487));
HA_X1 i_3446 (.CO (n_3728), .S (n_3727), .A (n_3515), .B (n_3508));
HA_X1 i_3442 (.CO (n_3723), .S (n_3722), .A (n_3536), .B (n_3529));
HA_X1 i_3366 (.CO (n_3646), .S (n_3645), .A (n_3473), .B (n_3642));
HA_X1 i_3362 (.CO (n_3641), .S (n_3640), .A (n_3468), .B (n_3632));
HA_X1 i_3358 (.CO (n_3636), .S (n_3635), .A (n_3622), .B (n_3463));
HA_X1 i_3354 (.CO (n_3631), .S (n_3630), .A (n_3617), .B (n_3612));
HA_X1 i_3350 (.CO (n_3626), .S (n_3625), .A (n_3448), .B (n_3607));
HA_X1 i_3346 (.CO (n_3621), .S (n_3620), .A (n_3438), .B (n_3602));
HA_X1 i_3342 (.CO (n_3616), .S (n_3615), .A (n_3582), .B (n_3577));
HA_X1 i_3338 (.CO (n_3611), .S (n_3610), .A (n_3428), .B (n_3592));
HA_X1 i_3334 (.CO (n_3606), .S (n_3605), .A (n_3408), .B (n_3572));
HA_X1 i_3330 (.CO (n_3601), .S (n_3600), .A (n_3423), .B (n_3418));
HA_X1 i_3326 (.CO (n_3596), .S (n_3595), .A (n_3567), .B (n_3562));
HA_X1 i_3322 (.CO (n_3591), .S (n_3590), .A (n_3486), .B (n_3477));
HA_X1 i_3318 (.CO (n_3586), .S (n_3585), .A (n_3507), .B (n_3500));
HA_X1 i_3314 (.CO (n_3581), .S (n_3580), .A (n_3528), .B (n_3521));
HA_X1 i_3310 (.CO (n_3576), .S (n_3575), .A (n_3549), .B (n_3542));
HA_X1 i_3306 (.CO (n_3571), .S (n_3570), .A (n_3398), .B (n_3393));
HA_X1 i_3302 (.CO (n_3566), .S (n_3565), .A (n_3328), .B (n_3321));
HA_X1 i_3298 (.CO (n_3561), .S (n_3560), .A (n_3349), .B (n_3342));
HA_X1 i_3294 (.CO (n_3556), .S (n_3555), .A (n_3370), .B (n_3363));
HA_X1 i_3214 (.CO (n_3475), .S (n_3474), .A (n_3308), .B (n_3471));
HA_X1 i_3210 (.CO (n_3470), .S (n_3469), .A (n_3303), .B (n_3461));
HA_X1 i_3206 (.CO (n_3465), .S (n_3464), .A (n_3456), .B (n_3451));
HA_X1 i_3202 (.CO (n_3460), .S (n_3459), .A (n_3288), .B (n_3446));
HA_X1 i_3198 (.CO (n_3455), .S (n_3454), .A (n_3426), .B (n_3283));
HA_X1 i_3194 (.CO (n_3450), .S (n_3449), .A (n_3278), .B (n_3436));
HA_X1 i_3190 (.CO (n_3445), .S (n_3444), .A (n_3421), .B (n_3416));
HA_X1 i_3186 (.CO (n_3440), .S (n_3439), .A (n_3273), .B (n_3268));
HA_X1 i_3182 (.CO (n_3435), .S (n_3434), .A (n_3253), .B (n_3248));
HA_X1 i_3178 (.CO (n_3430), .S (n_3429), .A (n_3391), .B (n_3383));
HA_X1 i_3174 (.CO (n_3425), .S (n_3424), .A (n_3243), .B (n_3401));
HA_X1 i_3170 (.CO (n_3420), .S (n_3419), .A (n_3327), .B (n_3320));
HA_X1 i_3166 (.CO (n_3415), .S (n_3414), .A (n_3348), .B (n_3341));
HA_X1 i_3162 (.CO (n_3410), .S (n_3409), .A (n_3369), .B (n_3362));
HA_X1 i_3158 (.CO (n_3405), .S (n_3404), .A (n_3233), .B (n_3228));
HA_X1 i_3154 (.CO (n_3400), .S (n_3399), .A (n_3164), .B (n_3157));
HA_X1 i_3150 (.CO (n_3395), .S (n_3394), .A (n_3185), .B (n_3178));
HA_X1 i_3146 (.CO (n_3390), .S (n_3389), .A (n_3206), .B (n_3199));
HA_X1 i_3067 (.CO (n_3310), .S (n_3309), .A (n_3151), .B (n_3306));
HA_X1 i_3063 (.CO (n_3305), .S (n_3304), .A (n_3146), .B (n_3296));
HA_X1 i_3059 (.CO (n_3300), .S (n_3299), .A (n_3286), .B (n_3291));
HA_X1 i_3055 (.CO (n_3295), .S (n_3294), .A (n_3131), .B (n_3136));
HA_X1 i_3051 (.CO (n_3290), .S (n_3289), .A (n_3266), .B (n_3126));
HA_X1 i_3047 (.CO (n_3285), .S (n_3284), .A (n_3261), .B (n_3121));
HA_X1 i_3043 (.CO (n_3280), .S (n_3279), .A (n_3256), .B (n_3251));
HA_X1 i_3039 (.CO (n_3275), .S (n_3274), .A (n_3241), .B (n_3116));
HA_X1 i_3035 (.CO (n_3270), .S (n_3269), .A (n_3101), .B (n_3096));
HA_X1 i_3031 (.CO (n_3265), .S (n_3264), .A (n_3231), .B (n_3226));
HA_X1 i_3027 (.CO (n_3260), .S (n_3259), .A (n_3156), .B (n_3086));
HA_X1 i_3023 (.CO (n_3255), .S (n_3254), .A (n_3177), .B (n_3170));
HA_X1 i_3019 (.CO (n_3250), .S (n_3249), .A (n_3198), .B (n_3191));
HA_X1 i_3015 (.CO (n_3245), .S (n_3244), .A (n_3219), .B (n_3212));
HA_X1 i_3011 (.CO (n_3240), .S (n_3239), .A (n_3081), .B (n_3076));
HA_X1 i_3007 (.CO (n_3235), .S (n_3234), .A (n_3018), .B (n_3011));
HA_X1 i_3003 (.CO (n_3230), .S (n_3229), .A (n_3039), .B (n_3032));
HA_X1 i_2999 (.CO (n_3225), .S (n_3224), .A (n_3060), .B (n_3053));
HA_X1 i_2928 (.CO (n_3153), .S (n_3152), .A (n_2998), .B (n_3149));
HA_X1 i_2924 (.CO (n_3148), .S (n_3147), .A (n_3139), .B (n_2993));
HA_X1 i_2920 (.CO (n_3143), .S (n_3142), .A (n_3129), .B (n_2988));
HA_X1 i_2916 (.CO (n_3138), .S (n_3137), .A (n_3119), .B (n_2983));
HA_X1 i_2912 (.CO (n_3133), .S (n_3132), .A (n_3109), .B (n_2973));
HA_X1 i_2908 (.CO (n_3128), .S (n_3127), .A (n_3094), .B (n_2968));
HA_X1 i_2904 (.CO (n_3123), .S (n_3122), .A (n_2958), .B (n_3104));
HA_X1 i_2900 (.CO (n_3118), .S (n_3117), .A (n_2943), .B (n_3089));
HA_X1 i_2896 (.CO (n_3113), .S (n_3112), .A (n_3074), .B (n_2953));
HA_X1 i_2892 (.CO (n_3108), .S (n_3107), .A (n_2938), .B (n_3084));
HA_X1 i_2888 (.CO (n_3103), .S (n_3102), .A (n_3017), .B (n_3010));
HA_X1 i_2884 (.CO (n_3098), .S (n_3097), .A (n_3038), .B (n_3031));
HA_X1 i_2880 (.CO (n_3093), .S (n_3092), .A (n_3059), .B (n_3052));
HA_X1 i_2876 (.CO (n_3088), .S (n_3087), .A (n_2928), .B (n_2919));
HA_X1 i_2872 (.CO (n_3083), .S (n_3082), .A (n_2863), .B (n_2856));
HA_X1 i_2868 (.CO (n_3078), .S (n_3077), .A (n_2884), .B (n_2877));
HA_X1 i_2864 (.CO (n_3073), .S (n_3072), .A (n_2905), .B (n_2898));
HA_X1 i_2792 (.CO (n_3000), .S (n_2999), .A (n_2850), .B (n_2996));
HA_X1 i_2788 (.CO (n_2995), .S (n_2994), .A (n_2986), .B (n_2845));
HA_X1 i_2784 (.CO (n_2990), .S (n_2989), .A (n_2976), .B (n_2840));
HA_X1 i_2780 (.CO (n_2985), .S (n_2984), .A (n_2966), .B (n_2971));
HA_X1 i_2776 (.CO (n_2980), .S (n_2979), .A (n_2961), .B (n_2956));
HA_X1 i_2772 (.CO (n_2975), .S (n_2974), .A (n_2946), .B (n_2941));
HA_X1 i_2768 (.CO (n_2970), .S (n_2969), .A (n_2820), .B (n_2815));
HA_X1 i_2764 (.CO (n_2965), .S (n_2964), .A (n_2795), .B (n_2810));
HA_X1 i_2760 (.CO (n_2960), .S (n_2959), .A (n_2918), .B (n_2805));
HA_X1 i_2756 (.CO (n_2955), .S (n_2954), .A (n_2790), .B (n_2931));
HA_X1 i_2752 (.CO (n_2950), .S (n_2949), .A (n_2869), .B (n_2862));
HA_X1 i_2748 (.CO (n_2945), .S (n_2944), .A (n_2890), .B (n_2883));
HA_X1 i_2744 (.CO (n_2940), .S (n_2939), .A (n_2911), .B (n_2904));
HA_X1 i_2740 (.CO (n_2935), .S (n_2934), .A (n_2716), .B (n_2785));
HA_X1 i_2736 (.CO (n_2930), .S (n_2929), .A (n_2737), .B (n_2730));
HA_X1 i_2732 (.CO (n_2925), .S (n_2924), .A (n_2758), .B (n_2751));
HA_X1 i_2660 (.CO (n_2852), .S (n_2851), .A (n_2710), .B (n_2848));
HA_X1 i_2656 (.CO (n_2847), .S (n_2846), .A (n_2838), .B (n_2705));
HA_X1 i_2652 (.CO (n_2842), .S (n_2841), .A (n_2828), .B (n_2700));
HA_X1 i_2648 (.CO (n_2837), .S (n_2836), .A (n_2690), .B (n_2823));
HA_X1 i_2644 (.CO (n_2832), .S (n_2831), .A (n_2685), .B (n_2818));
HA_X1 i_2640 (.CO (n_2827), .S (n_2826), .A (n_2808), .B (n_2803));
HA_X1 i_2636 (.CO (n_2822), .S (n_2821), .A (n_2793), .B (n_2680));
HA_X1 i_2632 (.CO (n_2817), .S (n_2816), .A (n_2670), .B (n_2665));
HA_X1 i_2628 (.CO (n_2812), .S (n_2811), .A (n_2788), .B (n_2783));
HA_X1 i_2624 (.CO (n_2807), .S (n_2806), .A (n_2722), .B (n_2715));
HA_X1 i_2620 (.CO (n_2802), .S (n_2801), .A (n_2743), .B (n_2736));
HA_X1 i_2616 (.CO (n_2797), .S (n_2796), .A (n_2764), .B (n_2757));
HA_X1 i_2612 (.CO (n_2792), .S (n_2791), .A (n_2645), .B (n_2635));
HA_X1 i_2608 (.CO (n_2787), .S (n_2786), .A (n_2587), .B (n_2580));
HA_X1 i_2604 (.CO (n_2782), .S (n_2781), .A (n_2608), .B (n_2601));
HA_X1 i_2600 (.CO (n_2777), .S (n_2776), .A (n_2629), .B (n_2622));
HA_X1 i_2536 (.CO (n_2712), .S (n_2711), .A (n_2574), .B (n_2576));
HA_X1 i_2532 (.CO (n_2707), .S (n_2706), .A (n_2569), .B (n_2698));
HA_X1 i_2528 (.CO (n_2702), .S (n_2701), .A (n_2564), .B (n_2688));
HA_X1 i_2524 (.CO (n_2697), .S (n_2696), .A (n_2554), .B (n_2683));
HA_X1 i_2520 (.CO (n_2692), .S (n_2691), .A (n_2549), .B (n_2678));
HA_X1 i_2516 (.CO (n_2687), .S (n_2686), .A (n_2668), .B (n_2663));
HA_X1 i_2512 (.CO (n_2682), .S (n_2681), .A (n_2653), .B (n_2544));
HA_X1 i_2508 (.CO (n_2677), .S (n_2676), .A (n_2534), .B (n_2529));
HA_X1 i_2504 (.CO (n_2672), .S (n_2671), .A (n_2579), .B (n_2648));
HA_X1 i_2500 (.CO (n_2667), .S (n_2666), .A (n_2600), .B (n_2593));
HA_X1 i_2496 (.CO (n_2662), .S (n_2661), .A (n_2621), .B (n_2614));
HA_X1 i_2492 (.CO (n_2657), .S (n_2656), .A (n_2505), .B (n_2634));
HA_X1 i_2488 (.CO (n_2652), .S (n_2651), .A (n_2449), .B (n_2519));
HA_X1 i_2484 (.CO (n_2647), .S (n_2646), .A (n_2470), .B (n_2463));
HA_X1 i_2480 (.CO (n_2642), .S (n_2641), .A (n_2491), .B (n_2484));
HA_X1 i_2415 (.CO (n_2576), .S (n_2575), .A (n_2443), .B (n_2572));
HA_X1 i_2411 (.CO (n_2571), .S (n_2570), .A (n_2562), .B (n_2438));
HA_X1 i_2407 (.CO (n_2566), .S (n_2565), .A (n_2433), .B (n_2552));
HA_X1 i_2403 (.CO (n_2561), .S (n_2560), .A (n_2542), .B (n_2423));
HA_X1 i_2399 (.CO (n_2556), .S (n_2555), .A (n_2537), .B (n_2418));
HA_X1 i_2395 (.CO (n_2551), .S (n_2550), .A (n_2413), .B (n_2532));
HA_X1 i_2391 (.CO (n_2546), .S (n_2545), .A (n_2403), .B (n_2398));
HA_X1 i_2387 (.CO (n_2541), .S (n_2540), .A (n_2512), .B (n_2504));
HA_X1 i_2383 (.CO (n_2536), .S (n_2535), .A (n_2448), .B (n_2393));
HA_X1 i_2379 (.CO (n_2531), .S (n_2530), .A (n_2469), .B (n_2462));
HA_X1 i_2375 (.CO (n_2526), .S (n_2525), .A (n_2490), .B (n_2483));
HA_X1 i_2371 (.CO (n_2521), .S (n_2520), .A (n_2388), .B (n_2383));
HA_X1 i_2367 (.CO (n_2516), .S (n_2515), .A (n_2340), .B (n_2333));
HA_X1 i_2363 (.CO (n_2511), .S (n_2510), .A (n_2361), .B (n_2354));
HA_X1 i_2298 (.CO (n_2445), .S (n_2444), .A (n_2320), .B (n_2441));
HA_X1 i_2294 (.CO (n_2440), .S (n_2439), .A (n_2431), .B (n_2315));
HA_X1 i_2290 (.CO (n_2435), .S (n_2434), .A (n_2421), .B (n_2310));
HA_X1 i_2286 (.CO (n_2430), .S (n_2429), .A (n_2416), .B (n_2411));
HA_X1 i_2282 (.CO (n_2425), .S (n_2424), .A (n_2401), .B (n_2396));
HA_X1 i_2278 (.CO (n_2420), .S (n_2419), .A (n_2295), .B (n_2290));
HA_X1 i_2274 (.CO (n_2415), .S (n_2414), .A (n_2280), .B (n_2275));
HA_X1 i_2270 (.CO (n_2410), .S (n_2409), .A (n_2386), .B (n_2381));
HA_X1 i_2266 (.CO (n_2405), .S (n_2404), .A (n_2339), .B (n_2332));
HA_X1 i_2262 (.CO (n_2400), .S (n_2399), .A (n_2360), .B (n_2353));
HA_X1 i_2258 (.CO (n_2395), .S (n_2394), .A (n_2255), .B (n_2374));
HA_X1 i_2254 (.CO (n_2390), .S (n_2389), .A (n_2207), .B (n_2270));
HA_X1 i_2250 (.CO (n_2385), .S (n_2384), .A (n_2228), .B (n_2221));
HA_X1 i_2246 (.CO (n_2380), .S (n_2379), .A (n_2249), .B (n_2242));
HA_X1 i_2189 (.CO (n_2322), .S (n_2321), .A (n_2201), .B (n_2318));
HA_X1 i_2185 (.CO (n_2317), .S (n_2316), .A (n_2308), .B (n_2196));
HA_X1 i_2181 (.CO (n_2312), .S (n_2311), .A (n_2298), .B (n_2191));
HA_X1 i_2177 (.CO (n_2307), .S (n_2306), .A (n_2181), .B (n_2293));
HA_X1 i_2173 (.CO (n_2302), .S (n_2301), .A (n_2283), .B (n_2278));
HA_X1 i_2169 (.CO (n_2297), .S (n_2296), .A (n_2273), .B (n_2176));
HA_X1 i_2165 (.CO (n_2292), .S (n_2291), .A (n_2263), .B (n_2166));
HA_X1 i_2161 (.CO (n_2287), .S (n_2286), .A (n_2206), .B (n_2156));
HA_X1 i_2157 (.CO (n_2282), .S (n_2281), .A (n_2227), .B (n_2220));
HA_X1 i_2153 (.CO (n_2277), .S (n_2276), .A (n_2248), .B (n_2241));
HA_X1 i_2149 (.CO (n_2272), .S (n_2271), .A (n_2151), .B (n_2142));
HA_X1 i_2145 (.CO (n_2267), .S (n_2266), .A (n_2107), .B (n_2100));
HA_X1 i_2141 (.CO (n_2262), .S (n_2261), .A (n_2128), .B (n_2121));
HA_X1 i_2083 (.CO (n_2203), .S (n_2202), .A (n_2087), .B (n_2199));
HA_X1 i_2079 (.CO (n_2198), .S (n_2197), .A (n_2082), .B (n_2189));
HA_X1 i_2075 (.CO (n_2193), .S (n_2192), .A (n_2072), .B (n_2077));
HA_X1 i_2071 (.CO (n_2188), .S (n_2187), .A (n_2067), .B (n_2179));
HA_X1 i_2067 (.CO (n_2183), .S (n_2182), .A (n_2169), .B (n_2164));
HA_X1 i_2063 (.CO (n_2178), .S (n_2177), .A (n_2052), .B (n_2047));
HA_X1 i_2059 (.CO (n_2173), .S (n_2172), .A (n_2149), .B (n_2141));
HA_X1 i_2055 (.CO (n_2168), .S (n_2167), .A (n_2099), .B (n_2092));
HA_X1 i_2051 (.CO (n_2163), .S (n_2162), .A (n_2120), .B (n_2113));
HA_X1 i_2047 (.CO (n_2158), .S (n_2157), .A (n_2037), .B (n_2134));
HA_X1 i_2043 (.CO (n_2153), .S (n_2152), .A (n_1994), .B (n_1987));
HA_X1 i_2039 (.CO (n_2148), .S (n_2147), .A (n_2015), .B (n_2008));
HA_X1 i_1981 (.CO (n_2089), .S (n_2088), .A (n_1981), .B (n_1983));
HA_X1 i_1977 (.CO (n_2084), .S (n_2083), .A (n_1976), .B (n_2075));
HA_X1 i_1973 (.CO (n_2079), .S (n_2078), .A (n_1966), .B (n_1971));
HA_X1 i_1969 (.CO (n_2074), .S (n_2073), .A (n_2050), .B (n_2065));
HA_X1 i_1965 (.CO (n_2069), .S (n_2068), .A (n_1961), .B (n_1956));
HA_X1 i_1961 (.CO (n_2064), .S (n_2063), .A (n_1951), .B (n_1946));
HA_X1 i_1957 (.CO (n_2059), .S (n_2058), .A (n_1941), .B (n_2040));
HA_X1 i_1953 (.CO (n_2054), .S (n_2053), .A (n_2000), .B (n_1993));
HA_X1 i_1949 (.CO (n_2049), .S (n_2048), .A (n_2021), .B (n_2014));
HA_X1 i_1945 (.CO (n_2044), .S (n_2043), .A (n_1936), .B (n_1926));
HA_X1 i_1941 (.CO (n_2039), .S (n_2038), .A (n_1899), .B (n_1892));
HA_X1 i_1937 (.CO (n_2034), .S (n_2033), .A (n_1920), .B (n_1913));
HA_X1 i_1887 (.CO (n_1983), .S (n_1982), .A (n_1879), .B (n_1979));
HA_X1 i_1883 (.CO (n_1978), .S (n_1977), .A (n_1969), .B (n_1874));
HA_X1 i_1879 (.CO (n_1973), .S (n_1972), .A (n_1959), .B (n_1869));
HA_X1 i_1875 (.CO (n_1968), .S (n_1967), .A (n_1949), .B (n_1944));
HA_X1 i_1871 (.CO (n_1963), .S (n_1962), .A (n_1854), .B (n_1859));
HA_X1 i_1867 (.CO (n_1958), .S (n_1957), .A (n_1934), .B (n_1849));
HA_X1 i_1863 (.CO (n_1953), .S (n_1952), .A (n_1891), .B (n_1884));
HA_X1 i_1859 (.CO (n_1948), .S (n_1947), .A (n_1912), .B (n_1905));
HA_X1 i_1855 (.CO (n_1943), .S (n_1942), .A (n_1830), .B (n_1925));
HA_X1 i_1851 (.CO (n_1938), .S (n_1937), .A (n_1795), .B (n_1788));
HA_X1 i_1847 (.CO (n_1933), .S (n_1932), .A (n_1816), .B (n_1809));
HA_X1 i_1796 (.CO (n_1881), .S (n_1880), .A (n_1782), .B (n_1877));
HA_X1 i_1792 (.CO (n_1876), .S (n_1875), .A (n_1777), .B (n_1867));
HA_X1 i_1788 (.CO (n_1871), .S (n_1870), .A (n_1857), .B (n_1772));
HA_X1 i_1784 (.CO (n_1866), .S (n_1865), .A (n_1762), .B (n_1852));
HA_X1 i_1780 (.CO (n_1861), .S (n_1860), .A (n_1752), .B (n_1842));
HA_X1 i_1776 (.CO (n_1856), .S (n_1855), .A (n_1837), .B (n_1829));
HA_X1 i_1772 (.CO (n_1851), .S (n_1850), .A (n_1794), .B (n_1787));
HA_X1 i_1768 (.CO (n_1846), .S (n_1845), .A (n_1815), .B (n_1808));
HA_X1 i_1764 (.CO (n_1841), .S (n_1840), .A (n_1699), .B (n_1742));
HA_X1 i_1760 (.CO (n_1836), .S (n_1835), .A (n_1720), .B (n_1713));
HA_X1 i_1709 (.CO (n_1784), .S (n_1783), .A (n_1693), .B (n_1695));
HA_X1 i_1705 (.CO (n_1779), .S (n_1778), .A (n_1688), .B (n_1770));
HA_X1 i_1701 (.CO (n_1774), .S (n_1773), .A (n_1760), .B (n_1765));
HA_X1 i_1697 (.CO (n_1769), .S (n_1768), .A (n_1678), .B (n_1755));
HA_X1 i_1693 (.CO (n_1764), .S (n_1763), .A (n_1740), .B (n_1673));
HA_X1 i_1689 (.CO (n_1759), .S (n_1758), .A (n_1698), .B (n_1663));
HA_X1 i_1685 (.CO (n_1754), .S (n_1753), .A (n_1719), .B (n_1712));
HA_X1 i_1681 (.CO (n_1749), .S (n_1748), .A (n_1648), .B (n_1733));
HA_X1 i_1677 (.CO (n_1744), .S (n_1743), .A (n_1621), .B (n_1614));
HA_X1 i_1673 (.CO (n_1739), .S (n_1738), .A (n_1642), .B (n_1635));
HA_X1 i_1630 (.CO (n_1695), .S (n_1694), .A (n_1608), .B (n_1610));
HA_X1 i_1626 (.CO (n_1690), .S (n_1689), .A (n_1681), .B (n_1603));
HA_X1 i_1622 (.CO (n_1685), .S (n_1684), .A (n_1666), .B (n_1676));
HA_X1 i_1618 (.CO (n_1680), .S (n_1679), .A (n_1661), .B (n_1593));
HA_X1 i_1614 (.CO (n_1675), .S (n_1674), .A (n_1656), .B (n_1588));
HA_X1 i_1610 (.CO (n_1670), .S (n_1669), .A (n_1627), .B (n_1620));
HA_X1 i_1606 (.CO (n_1665), .S (n_1664), .A (n_1647), .B (n_1641));
HA_X1 i_1602 (.CO (n_1660), .S (n_1659), .A (n_1534), .B (n_1578));
HA_X1 i_1598 (.CO (n_1655), .S (n_1654), .A (n_1555), .B (n_1548));
HA_X1 i_1554 (.CO (n_1610), .S (n_1609), .A (n_1528), .B (n_1530));
HA_X1 i_1550 (.CO (n_1605), .S (n_1604), .A (n_1523), .B (n_1596));
HA_X1 i_1546 (.CO (n_1600), .S (n_1599), .A (n_1581), .B (n_1518));
HA_X1 i_1542 (.CO (n_1595), .S (n_1594), .A (n_1508), .B (n_1513));
HA_X1 i_1538 (.CO (n_1590), .S (n_1589), .A (n_1503), .B (n_1576));
HA_X1 i_1534 (.CO (n_1585), .S (n_1584), .A (n_1547), .B (n_1540));
HA_X1 i_1530 (.CO (n_1580), .S (n_1579), .A (n_1498), .B (n_1561));
HA_X1 i_1526 (.CO (n_1575), .S (n_1574), .A (n_1476), .B (n_1469));
HA_X1 i_1482 (.CO (n_1530), .S (n_1529), .A (n_1456), .B (n_1458));
HA_X1 i_1478 (.CO (n_1525), .S (n_1524), .A (n_1516), .B (n_1451));
HA_X1 i_1474 (.CO (n_1520), .S (n_1519), .A (n_1446), .B (n_1511));
HA_X1 i_1470 (.CO (n_1515), .S (n_1514), .A (n_1441), .B (n_1436));
HA_X1 i_1466 (.CO (n_1510), .S (n_1509), .A (n_1468), .B (n_1461));
HA_X1 i_1462 (.CO (n_1505), .S (n_1504), .A (n_1489), .B (n_1482));
HA_X1 i_1458 (.CO (n_1500), .S (n_1499), .A (n_1394), .B (n_1431));
HA_X1 i_1454 (.CO (n_1495), .S (n_1494), .A (n_1415), .B (n_1408));
HA_X1 i_1418 (.CO (n_1458), .S (n_1457), .A (n_1449), .B (n_1390));
HA_X1 i_1414 (.CO (n_1453), .S (n_1452), .A (n_1444), .B (n_1383));
HA_X1 i_1410 (.CO (n_1448), .S (n_1447), .A (n_1378), .B (n_1439));
HA_X1 i_1406 (.CO (n_1443), .S (n_1442), .A (n_1368), .B (n_1429));
HA_X1 i_1402 (.CO (n_1438), .S (n_1437), .A (n_1407), .B (n_1400));
HA_X1 i_1398 (.CO (n_1433), .S (n_1432), .A (n_1359), .B (n_1420));
HA_X1 i_1394 (.CO (n_1428), .S (n_1427), .A (n_1345), .B (n_1338));
HA_X1 i_1357 (.CO (n_1390), .S (n_1389), .A (n_1325), .B (n_1327));
HA_X1 i_1353 (.CO (n_1385), .S (n_1384), .A (n_1320), .B (n_1376));
HA_X1 i_1349 (.CO (n_1380), .S (n_1379), .A (n_1310), .B (n_1315));
HA_X1 i_1345 (.CO (n_1375), .S (n_1374), .A (n_1330), .B (n_1366));
HA_X1 i_1341 (.CO (n_1370), .S (n_1369), .A (n_1351), .B (n_1344));
HA_X1 i_1337 (.CO (n_1365), .S (n_1364), .A (n_1283), .B (n_1276));
HA_X1 i_1300 (.CO (n_1327), .S (n_1326), .A (n_1272), .B (n_1270));
HA_X1 i_1296 (.CO (n_1322), .S (n_1321), .A (n_1313), .B (n_1308));
HA_X1 i_1292 (.CO (n_1317), .S (n_1316), .A (n_1303), .B (n_1260));
HA_X1 i_1288 (.CO (n_1312), .S (n_1311), .A (n_1282), .B (n_1275));
HA_X1 i_1284 (.CO (n_1307), .S (n_1306), .A (n_1245), .B (n_1296));
HA_X1 i_1280 (.CO (n_1302), .S (n_1301), .A (n_1239), .B (n_1232));
HA_X1 i_1251 (.CO (n_1272), .S (n_1271), .A (n_1221), .B (n_1219));
HA_X1 i_1247 (.CO (n_1267), .S (n_1266), .A (n_1214), .B (n_1258));
HA_X1 i_1243 (.CO (n_1262), .S (n_1261), .A (n_1224), .B (n_1253));
HA_X1 i_1239 (.CO (n_1257), .S (n_1256), .A (n_1244), .B (n_1238));
HA_X1 i_1235 (.CO (n_1252), .S (n_1251), .A (n_1186), .B (n_1179));
HA_X1 i_1205 (.CO (n_1221), .S (n_1220), .A (n_1175), .B (n_1173));
HA_X1 i_1201 (.CO (n_1216), .S (n_1215), .A (n_1168), .B (n_1207));
HA_X1 i_1197 (.CO (n_1211), .S (n_1210), .A (n_1178), .B (n_1163));
HA_X1 i_1193 (.CO (n_1206), .S (n_1205), .A (n_1141), .B (n_1192));
HA_X1 i_1163 (.CO (n_1175), .S (n_1174), .A (n_1135), .B (n_1166));
HA_X1 i_1159 (.CO (n_1170), .S (n_1169), .A (n_1161), .B (n_1130));
HA_X1 i_1155 (.CO (n_1165), .S (n_1164), .A (n_1154), .B (n_1147));
HA_X1 i_1151 (.CO (n_1160), .S (n_1159), .A (n_1114), .B (n_1107));
HA_X1 i_1129 (.CO (n_1137), .S (n_1136), .A (n_1128), .B (n_1101));
HA_X1 i_1125 (.CO (n_1132), .S (n_1131), .A (n_1113), .B (n_1106));
HA_X1 i_1121 (.CO (n_1127), .S (n_1126), .A (n_1078), .B (n_1092));
HA_X1 i_1098 (.CO (n_1103), .S (n_1102), .A (n_1074), .B (n_1072));
HA_X1 i_1094 (.CO (n_1098), .S (n_1097), .A (n_1084), .B (n_1077));
HA_X1 i_1071 (.CO (n_1074), .S (n_1073), .A (n_1056), .B (n_1053));
HA_X1 i_1067 (.CO (n_1069), .S (n_1068), .A (n_1040), .B (n_1046));
HA_X1 i_1052 (.CO (n_1053), .S (n_1052), .A (n_1030), .B (n_1045));

endmodule //datapath

module multiplyTimes (inputA, inputB, result);

output [63:0] result;
input [31:0] inputA;
input [31:0] inputB;


datapath i_0 (.result ({result[63], result[62], result[61], result[60], result[59], 
    result[58], result[57], result[56], result[55], result[54], result[53], result[52], 
    result[51], result[50], result[49], result[48], result[47], result[46], result[45], 
    result[44], result[43], result[42], result[41], result[40], result[39], result[38], 
    result[37], result[36], result[35], result[34], result[33], result[32], result[31], 
    result[30], result[29], result[28], result[27], result[26], result[25], result[24], 
    result[23], result[22], result[21], result[20], result[19], result[18], result[17], 
    result[16], result[15], result[14], result[13], result[12], result[11], result[10], 
    result[9], result[8], result[7], result[6], result[5], result[4], result[3], 
    result[2], result[1], result[0]}), .inputA ({inputA[31], inputA[30], inputA[29], 
    inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], inputA[22], 
    inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], inputA[15], 
    inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], inputA[8], 
    inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], inputA[1], 
    inputA[0]}), .inputB ({inputB[31], inputB[30], inputB[29], inputB[28], inputB[27], 
    inputB[26], inputB[25], inputB[24], inputB[23], inputB[22], inputB[21], inputB[20], 
    inputB[19], inputB[18], inputB[17], inputB[16], inputB[15], inputB[14], inputB[13], 
    inputB[12], inputB[11], inputB[10], inputB[9], inputB[8], inputB[7], inputB[6], 
    inputB[5], inputB[4], inputB[3], inputB[2], inputB[1], inputB[0]}));

endmodule //multiplyTimes

module integrationMult (clk, reset, en, inputA, inputB, result);

output [63:0] result;
input clk;
input en;
input [31:0] inputA;
input [31:0] inputB;
input reset;
wire CTS_n3;
wire \outB_reg[31] ;
wire \outB_reg[30] ;
wire \outB_reg[29] ;
wire \outB_reg[28] ;
wire \outB_reg[27] ;
wire \outB_reg[26] ;
wire \outB_reg[25] ;
wire \outB_reg[24] ;
wire \outB_reg[23] ;
wire \outB_reg[22] ;
wire \outB_reg[21] ;
wire \outB_reg[20] ;
wire \outB_reg[19] ;
wire \outB_reg[18] ;
wire \outB_reg[17] ;
wire \outB_reg[16] ;
wire \outB_reg[15] ;
wire \outB_reg[14] ;
wire \outB_reg[13] ;
wire \outB_reg[12] ;
wire \outB_reg[11] ;
wire \outB_reg[10] ;
wire \outB_reg[9] ;
wire \outB_reg[8] ;
wire \outB_reg[7] ;
wire \outB_reg[6] ;
wire \outB_reg[5] ;
wire \outB_reg[4] ;
wire \outB_reg[3] ;
wire \outB_reg[2] ;
wire \outB_reg[1] ;
wire \outB_reg[0] ;
wire \outA_reg[31] ;
wire \outA_reg[30] ;
wire \outA_reg[29] ;
wire \outA_reg[28] ;
wire \outA_reg[27] ;
wire \outA_reg[26] ;
wire \outA_reg[25] ;
wire \outA_reg[24] ;
wire \outA_reg[23] ;
wire \outA_reg[22] ;
wire \outA_reg[21] ;
wire \outA_reg[20] ;
wire \outA_reg[19] ;
wire \outA_reg[18] ;
wire \outA_reg[17] ;
wire \outA_reg[16] ;
wire \outA_reg[15] ;
wire \outA_reg[14] ;
wire \outA_reg[13] ;
wire \outA_reg[12] ;
wire \outA_reg[11] ;
wire \outA_reg[10] ;
wire \outA_reg[9] ;
wire \outA_reg[8] ;
wire \outA_reg[7] ;
wire \outA_reg[6] ;
wire \outA_reg[5] ;
wire \outA_reg[4] ;
wire \outA_reg[3] ;
wire \outA_reg[2] ;
wire \outA_reg[1] ;
wire \outA_reg[0] ;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;


registerNbits outA (.out ({result[31], result[30], result[29], result[28], result[27], 
    result[26], result[25], result[24], result[23], result[22], result[21], result[20], 
    result[19], result[18], result[17], result[16], result[15], result[14], result[13], 
    result[12], result[11], result[10], result[9], result[8], result[7], result[6], 
    result[5], result[4], result[3], result[2], result[1], result[0]}), .en (en), .inp ({
    \outB_reg[31] , \outB_reg[30] , \outB_reg[29] , \outB_reg[28] , \outB_reg[27] , 
    \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , \outB_reg[23] , \outB_reg[22] , 
    \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , \outB_reg[18] , \outB_reg[17] , 
    \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , \outB_reg[13] , \outB_reg[12] , 
    \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , \outB_reg[8] , \outB_reg[7] , 
    \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , 
    \outB_reg[0] }), .reset (reset), .clk_CTSPP_2 (clk));
registerNbits__2_8 outB (.out ({result[63], result[62], result[61], result[60], result[59], 
    result[58], result[57], result[56], result[55], result[54], result[53], result[52], 
    result[51], result[50], result[49], result[48], result[47], result[46], result[45], 
    result[44], result[43], result[42], result[41], result[40], result[39], result[38], 
    result[37], result[36], result[35], result[34], result[33], result[32]}), .clk_CTSPP_0 (CTS_n3)
    , .en (en), .inp ({\outA_reg[31] , \outA_reg[30] , \outA_reg[29] , \outA_reg[28] , 
    \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , \outA_reg[24] , \outA_reg[23] , 
    \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , \outA_reg[19] , \outA_reg[18] , 
    \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , \outA_reg[14] , \outA_reg[13] , 
    \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , \outA_reg[9] , \outA_reg[8] , 
    \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , 
    \outA_reg[1] , \outA_reg[0] }), .reset (reset), .clk_CTSPP_2 (clk));
registerNbits__2_5 regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , 
    \B_reg[27] , \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , 
    \B_reg[21] , \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , 
    \B_reg[15] , \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , 
    \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .en (en), .inp ({inputB[31], inputB[30], 
    inputB[29], inputB[28], inputB[27], inputB[26], inputB[25], inputB[24], inputB[23], 
    inputB[22], inputB[21], inputB[20], inputB[19], inputB[18], inputB[17], inputB[16], 
    inputB[15], inputB[14], inputB[13], inputB[12], inputB[11], inputB[10], inputB[9], 
    inputB[8], inputB[7], inputB[6], inputB[5], inputB[4], inputB[3], inputB[2], 
    inputB[1], inputB[0]}), .reset (reset), .clk_CTSPP_0 (CTS_n3));
registerNbits__2_2 regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .en (en), .inp ({inputA[31], inputA[30], 
    inputA[29], inputA[28], inputA[27], inputA[26], inputA[25], inputA[24], inputA[23], 
    inputA[22], inputA[21], inputA[20], inputA[19], inputA[18], inputA[17], inputA[16], 
    inputA[15], inputA[14], inputA[13], inputA[12], inputA[11], inputA[10], inputA[9], 
    inputA[8], inputA[7], inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], 
    inputA[1], inputA[0]}), .reset (reset), .clk_CTSPP_0 (CTS_n3));
multiplyTimes mult (.result ({\outA_reg[31] , \outA_reg[30] , \outA_reg[29] , \outA_reg[28] , 
    \outA_reg[27] , \outA_reg[26] , \outA_reg[25] , \outA_reg[24] , \outA_reg[23] , 
    \outA_reg[22] , \outA_reg[21] , \outA_reg[20] , \outA_reg[19] , \outA_reg[18] , 
    \outA_reg[17] , \outA_reg[16] , \outA_reg[15] , \outA_reg[14] , \outA_reg[13] , 
    \outA_reg[12] , \outA_reg[11] , \outA_reg[10] , \outA_reg[9] , \outA_reg[8] , 
    \outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , 
    \outA_reg[1] , \outA_reg[0] , \outB_reg[31] , \outB_reg[30] , \outB_reg[29] , 
    \outB_reg[28] , \outB_reg[27] , \outB_reg[26] , \outB_reg[25] , \outB_reg[24] , 
    \outB_reg[23] , \outB_reg[22] , \outB_reg[21] , \outB_reg[20] , \outB_reg[19] , 
    \outB_reg[18] , \outB_reg[17] , \outB_reg[16] , \outB_reg[15] , \outB_reg[14] , 
    \outB_reg[13] , \outB_reg[12] , \outB_reg[11] , \outB_reg[10] , \outB_reg[9] , 
    \outB_reg[8] , \outB_reg[7] , \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , 
    \outB_reg[2] , \outB_reg[1] , \outB_reg[0] }), .inputA ({\A_reg[31] , \A_reg[30] , 
    \A_reg[29] , \A_reg[28] , \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , 
    \A_reg[23] , \A_reg[22] , \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , 
    \A_reg[17] , \A_reg[16] , \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , 
    \A_reg[11] , \A_reg[10] , \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , 
    \A_reg[4] , \A_reg[3] , \A_reg[2] , \A_reg[1] , \A_reg[0] }), .inputB ({\B_reg[31] , 
    \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , \B_reg[26] , \B_reg[25] , 
    \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , \B_reg[20] , \B_reg[19] , 
    \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , \B_reg[14] , \B_reg[13] , 
    \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , \B_reg[8] , \B_reg[7] , \B_reg[6] , 
    \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] }));

endmodule //integrationMult


