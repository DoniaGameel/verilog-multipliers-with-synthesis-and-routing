
// 	Wed Jan  4 02:22:52 2023
//	vlsi
//	localhost.localdomain

module datapath__0_4 (p_0, p_1, MP_final);

output [22:0] MP_final;
input [22:0] p_0;
input [22:0] p_1;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;


AND2_X1 i_44 (.ZN (n_21), .A1 (n_12), .A2 (p_1[13]));
AND2_X1 i_43 (.ZN (n_20), .A1 (p_1[14]), .A2 (n_21));
AND2_X1 i_41 (.ZN (n_19), .A1 (p_1[15]), .A2 (n_20));
AND2_X1 i_39 (.ZN (n_18), .A1 (p_1[16]), .A2 (n_19));
AND2_X1 i_37 (.ZN (n_17), .A1 (p_1[17]), .A2 (n_18));
AND2_X1 i_35 (.ZN (n_16), .A1 (p_1[18]), .A2 (n_17));
AND2_X1 i_33 (.ZN (n_15), .A1 (p_1[19]), .A2 (n_16));
AND2_X1 i_31 (.ZN (n_14), .A1 (p_1[20]), .A2 (n_15));
NAND2_X1 i_29 (.ZN (n_13), .A1 (p_1[21]), .A2 (n_14));
XNOR2_X1 i_27 (.ZN (MP_final[22]), .A (p_1[22]), .B (n_13));
XOR2_X1 i_42 (.Z (MP_final[21]), .A (p_1[21]), .B (n_14));
XOR2_X1 i_40 (.Z (MP_final[20]), .A (p_1[20]), .B (n_15));
XOR2_X1 i_38 (.Z (MP_final[19]), .A (p_1[19]), .B (n_16));
XOR2_X1 i_36 (.Z (MP_final[18]), .A (p_1[18]), .B (n_17));
XOR2_X1 i_34 (.Z (MP_final[17]), .A (p_1[17]), .B (n_18));
XOR2_X1 i_32 (.Z (MP_final[16]), .A (p_1[16]), .B (n_19));
XOR2_X1 i_30 (.Z (MP_final[15]), .A (p_1[15]), .B (n_20));
XOR2_X1 i_28 (.Z (MP_final[14]), .A (p_1[14]), .B (n_21));
XOR2_X1 i_26 (.Z (MP_final[13]), .A (p_1[13]), .B (n_12));
AND2_X1 i_25 (.ZN (n_12), .A1 (n_11), .A2 (p_1[12]));
XOR2_X1 i_24 (.Z (MP_final[12]), .A (p_1[12]), .B (n_11));
AND2_X1 i_23 (.ZN (n_11), .A1 (n_10), .A2 (p_1[11]));
XOR2_X1 i_22 (.Z (MP_final[11]), .A (p_1[11]), .B (n_10));
AND2_X1 i_21 (.ZN (n_10), .A1 (n_9), .A2 (p_1[10]));
XOR2_X1 i_20 (.Z (MP_final[10]), .A (p_1[10]), .B (n_9));
AND2_X1 i_19 (.ZN (n_9), .A1 (n_8), .A2 (p_1[9]));
XOR2_X1 i_18 (.Z (MP_final[9]), .A (p_1[9]), .B (n_8));
AND2_X1 i_17 (.ZN (n_8), .A1 (n_7), .A2 (p_1[8]));
XOR2_X1 i_16 (.Z (MP_final[8]), .A (p_1[8]), .B (n_7));
AND2_X1 i_15 (.ZN (n_7), .A1 (n_6), .A2 (p_1[7]));
XOR2_X1 i_14 (.Z (MP_final[7]), .A (p_1[7]), .B (n_6));
AND2_X1 i_13 (.ZN (n_6), .A1 (n_5), .A2 (p_1[6]));
XOR2_X1 i_12 (.Z (MP_final[6]), .A (p_1[6]), .B (n_5));
AND2_X1 i_11 (.ZN (n_5), .A1 (n_4), .A2 (p_1[5]));
XOR2_X1 i_10 (.Z (MP_final[5]), .A (p_1[5]), .B (n_4));
AND2_X1 i_9 (.ZN (n_4), .A1 (n_3), .A2 (p_1[4]));
XOR2_X1 i_8 (.Z (MP_final[4]), .A (p_1[4]), .B (n_3));
AND2_X1 i_7 (.ZN (n_3), .A1 (n_2), .A2 (p_1[3]));
XOR2_X1 i_6 (.Z (MP_final[3]), .A (p_1[3]), .B (n_2));
AND2_X1 i_5 (.ZN (n_2), .A1 (n_1), .A2 (p_1[2]));
XOR2_X1 i_4 (.Z (MP_final[2]), .A (p_1[2]), .B (n_1));
AND2_X1 i_3 (.ZN (n_1), .A1 (n_0), .A2 (p_1[1]));
XOR2_X1 i_2 (.Z (MP_final[1]), .A (p_1[1]), .B (n_0));
AND2_X1 i_1 (.ZN (n_0), .A1 (p_1[0]), .A2 (p_0[0]));
XOR2_X1 i_0 (.Z (MP_final[0]), .A (p_0[0]), .B (p_1[0]));

endmodule //datapath__0_4

module Reg (in, clk, out);

output [31:0] out;
input clk;
input [31:0] in;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk), .D (in[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk), .D (in[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk), .D (in[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk), .D (in[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk), .D (in[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk), .D (in[11]));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (clk), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk), .D (in[13]));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (clk), .D (in[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk), .D (in[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk), .D (in[16]));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (clk), .D (in[17]));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (clk), .D (in[18]));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (clk), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk), .D (in[20]));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (clk), .D (in[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk), .D (in[31]));

endmodule //Reg

module datapath (B, A, Out);

output [47:0] Out;
input [23:0] A;
input [23:0] B;
wire n_20;
wire n_3;
wire n_19;
wire n_30;
wire n_1534;
wire n_29;
wire n_32;
wire n_424;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_25;
wire n_107;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_66;
wire n_150;
wire n_64;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_143;
wire n_141;
wire n_149;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_28;
wire n_170;
wire n_65;
wire n_99;
wire n_423;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_100;
wire n_421;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_386;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_422;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_417;
wire n_416;
wire n_144;
wire n_145;
wire n_393;
wire n_392;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_381;
wire n_380;
wire n_172;
wire n_173;
wire n_397;
wire n_391;
wire n_179;
wire n_180;
wire n_183;
wire n_454;
wire n_184;
wire n_185;
wire n_186;
wire n_388;
wire n_387;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_455;
wire n_331;
wire n_199;
wire n_200;
wire n_201;
wire n_340;
wire n_202;
wire n_203;
wire n_446;
wire n_445;
wire n_210;
wire n_211;
wire n_213;
wire n_370;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_223;
wire n_374;
wire n_224;
wire n_385;
wire n_225;
wire n_376;
wire n_390;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_1955;
wire n_389;
wire n_169;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_439;
wire n_437;
wire n_271;
wire n_375;
wire n_355;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_198;
wire n_299;
wire n_373;
wire n_371;
wire n_300;
wire n_369;
wire n_359;
wire n_358;
wire n_301;
wire n_302;
wire n_303;
wire n_321;
wire n_269;
wire n_310;
wire n_207;
wire n_208;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_427;
wire n_354;
wire n_322;
wire n_262;
wire n_263;
wire n_329;
wire n_174;
wire n_168;
wire n_171;
wire n_336;
wire n_337;
wire n_177;
wire n_178;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_189;
wire n_212;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_312;
wire n_305;
wire n_383;
wire n_276;
wire n_275;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_273;
wire n_268;
wire n_428;
wire n_429;
wire n_430;
wire n_309;
wire n_307;
wire n_306;
wire n_431;
wire n_281;
wire n_283;
wire n_270;
wire n_432;
wire n_433;
wire n_286;
wire n_434;
wire n_285;
wire n_284;
wire n_435;
wire n_436;
wire n_520;
wire n_523;
wire n_440;
wire n_517;
wire n_443;
wire n_534;
wire n_537;
wire n_447;
wire n_287;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_492;
wire n_489;
wire n_456;
wire n_466;
wire n_465;
wire n_463;
wire n_464;
wire n_541;
wire n_540;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_578;
wire n_490;
wire n_580;
wire n_491;
wire n_579;
wire n_493;
wire n_571;
wire n_568;
wire n_497;
wire n_569;
wire n_499;
wire n_500;
wire n_503;
wire n_502;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_304;
wire n_511;
wire n_274;
wire n_512;
wire n_513;
wire n_514;
wire n_614;
wire n_615;
wire n_518;
wire n_519;
wire n_565;
wire n_566;
wire n_525;
wire n_526;
wire n_527;
wire n_222;
wire n_528;
wire n_246;
wire n_267;
wire n_245;
wire n_529;
wire n_524;
wire n_516;
wire n_538;
wire n_539;
wire n_470;
wire n_462;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_495;
wire n_461;
wire n_563;
wire n_772;
wire n_773;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_576;
wire n_581;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_781;
wire n_782;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_556;
wire n_426;
wire n_639;
wire n_2243;
wire n_458;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_1339;
wire n_646;
wire n_1235;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_599;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_666;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_611;
wire n_460;
wire n_688;
wire n_777;
wire n_783;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_582;
wire n_713;
wire n_598;
wire n_714;
wire n_605;
wire n_604;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_560;
wire n_720;
wire n_721;
wire n_722;
wire n_607;
wire n_723;
wire n_724;
wire n_725;
wire n_31;
wire n_1532;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_1116;
wire n_732;
wire n_425;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_738;
wire n_1128;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_459;
wire n_606;
wire n_610;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_849;
wire n_848;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_802;
wire n_831;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_803;
wire n_913;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_1676;
wire n_818;
wire n_819;
wire n_820;
wire n_750;
wire n_821;
wire n_694;
wire n_761;
wire n_760;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_1120;
wire n_1017;
wire n_854;
wire n_1115;
wire n_1114;
wire n_858;
wire n_859;
wire n_1008;
wire n_861;
wire n_862;
wire n_863;
wire n_229;
wire n_864;
wire n_865;
wire n_866;
wire n_833;
wire n_867;
wire n_868;
wire n_832;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_843;
wire n_846;
wire n_844;
wire n_882;
wire n_883;
wire n_990;
wire n_989;
wire n_890;
wire n_891;
wire n_840;
wire n_834;
wire n_847;
wire n_841;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_1013;
wire n_1011;
wire n_900;
wire n_995;
wire n_994;
wire n_907;
wire n_908;
wire n_1022;
wire n_1021;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_1117;
wire n_1113;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_924;
wire n_906;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_912;
wire n_976;
wire n_909;
wire n_977;
wire n_928;
wire n_1232;
wire n_939;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_901;
wire n_997;
wire n_1052;
wire n_1010;
wire n_1053;
wire n_1012;
wire n_1035;
wire n_1019;
wire n_1020;
wire n_1103;
wire n_1097;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_940;
wire n_905;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1032;
wire n_1096;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_887;
wire n_899;
wire n_1123;
wire n_903;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1530;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1050;
wire n_1048;
wire n_1036;
wire n_1137;
wire n_884;
wire n_860;
wire n_855;
wire n_1138;
wire n_1139;
wire n_896;
wire n_902;
wire n_888;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1301;
wire n_1300;
wire n_1149;
wire n_1296;
wire n_1295;
wire n_1155;
wire n_1156;
wire n_1289;
wire n_1173;
wire n_1162;
wire n_1163;
wire n_1051;
wire n_1231;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1060;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_889;
wire n_1209;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1200;
wire n_1199;
wire n_1195;
wire n_1226;
wire n_1225;
wire n_1201;
wire n_1202;
wire n_1260;
wire n_1259;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1031;
wire n_1210;
wire n_904;
wire n_944;
wire n_1211;
wire n_1329;
wire n_1327;
wire n_1215;
wire n_949;
wire n_1216;
wire n_948;
wire n_1217;
wire n_947;
wire n_950;
wire n_1218;
wire n_1219;
wire n_1192;
wire n_1191;
wire n_1223;
wire n_1224;
wire n_1158;
wire n_1157;
wire n_1229;
wire n_1150;
wire n_1148;
wire n_1233;
wire n_1234;
wire n_1221;
wire n_1237;
wire n_1220;
wire n_1238;
wire n_1214;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_999;
wire n_1249;
wire n_955;
wire n_945;
wire n_978;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1061;
wire n_1056;
wire n_1063;
wire n_1062;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1292;
wire n_1264;
wire n_1265;
wire n_1711;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1144;
wire n_1304;
wire n_1306;
wire n_1030;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1418;
wire n_1420;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1479;
wire n_1481;
wire n_1340;
wire n_1478;
wire n_1342;
wire n_1484;
wire n_1485;
wire n_1347;
wire n_1482;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1441;
wire n_1426;
wire n_1436;
wire n_1379;
wire n_1380;
wire n_1385;
wire n_1236;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1239;
wire n_1400;
wire n_1263;
wire n_1401;
wire n_1362;
wire n_1365;
wire n_1407;
wire n_1408;
wire n_1501;
wire n_1461;
wire n_1416;
wire n_1417;
wire n_1423;
wire n_1442;
wire n_1427;
wire n_1428;
wire n_1429;
wire n_1430;
wire n_1431;
wire n_1432;
wire n_1375;
wire n_1433;
wire n_1434;
wire n_1435;
wire n_1344;
wire n_1631;
wire n_1437;
wire n_1438;
wire n_1439;
wire n_1440;
wire n_1526;
wire n_1341;
wire n_1445;
wire n_1446;
wire n_1371;
wire n_1372;
wire n_1451;
wire n_1505;
wire n_1504;
wire n_1457;
wire n_1458;
wire n_1462;
wire n_1522;
wire n_1463;
wire n_1464;
wire n_1465;
wire n_1466;
wire n_1467;
wire n_1468;
wire n_1469;
wire n_1470;
wire n_1471;
wire n_1472;
wire n_1473;
wire n_1474;
wire n_1196;
wire n_1145;
wire n_1475;
wire n_1326;
wire n_1338;
wire n_1486;
wire n_1487;
wire n_1488;
wire n_1489;
wire n_1490;
wire n_1491;
wire n_1492;
wire n_1493;
wire n_1494;
wire n_1495;
wire n_1496;
wire n_1497;
wire n_1498;
wire n_1499;
wire n_1500;
wire n_1413;
wire n_1443;
wire n_1510;
wire n_1511;
wire n_1512;
wire n_1513;
wire n_1514;
wire n_1515;
wire n_1516;
wire n_1517;
wire n_1518;
wire n_1519;
wire n_1520;
wire n_1502;
wire n_1450;
wire n_1536;
wire n_1537;
wire n_1538;
wire n_1319;
wire n_1321;
wire n_1323;
wire n_1539;
wire n_1540;
wire n_1541;
wire n_1542;
wire n_1543;
wire n_1544;
wire n_1545;
wire n_1546;
wire n_1547;
wire n_1548;
wire n_1549;
wire n_1550;
wire n_1551;
wire n_1552;
wire n_1616;
wire n_1615;
wire n_1556;
wire n_1601;
wire n_1604;
wire n_1602;
wire n_1564;
wire n_1565;
wire n_1587;
wire n_1508;
wire n_1570;
wire n_1571;
wire n_1572;
wire n_1636;
wire n_1635;
wire n_1578;
wire n_1786;
wire n_1581;
wire n_1029;
wire n_1317;
wire n_1792;
wire n_1582;
wire n_1583;
wire n_1318;
wire n_1584;
wire n_1585;
wire n_1627;
wire n_1626;
wire n_1591;
wire n_1592;
wire n_1593;
wire n_1594;
wire n_1595;
wire n_1596;
wire n_1597;
wire n_1598;
wire n_1599;
wire n_1600;
wire n_1655;
wire n_1658;
wire n_1618;
wire n_1619;
wire n_1731;
wire n_1710;
wire n_1625;
wire n_1745;
wire n_1746;
wire n_1791;
wire n_1632;
wire n_1633;
wire n_1612;
wire n_1611;
wire n_1637;
wire n_1638;
wire n_1639;
wire n_1449;
wire n_1641;
wire n_1642;
wire n_1643;
wire n_1644;
wire n_1645;
wire n_1646;
wire n_1788;
wire n_1787;
wire n_1651;
wire n_1762;
wire n_1648;
wire n_1656;
wire n_1657;
wire n_1739;
wire n_1738;
wire n_1663;
wire n_1664;
wire n_1665;
wire n_1666;
wire n_1444;
wire n_1667;
wire n_1509;
wire n_1503;
wire n_1521;
wire n_1525;
wire n_1668;
wire n_1669;
wire n_1670;
wire n_1671;
wire n_1672;
wire n_1673;
wire n_1674;
wire n_1675;
wire n_1881;
wire n_1677;
wire n_1678;
wire n_1679;
wire n_1680;
wire n_1681;
wire n_1682;
wire n_1683;
wire n_1684;
wire n_1685;
wire n_1686;
wire n_1687;
wire n_1688;
wire n_1689;
wire n_1690;
wire n_1691;
wire n_1692;
wire n_1693;
wire n_1694;
wire n_1695;
wire n_1696;
wire n_1697;
wire n_1662;
wire n_1717;
wire n_1727;
wire n_1448;
wire n_1729;
wire n_1734;
wire n_1730;
wire n_1735;
wire n_1825;
wire n_1573;
wire n_1741;
wire n_1742;
wire n_1784;
wire n_1760;
wire n_1747;
wire n_1748;
wire n_1749;
wire n_1750;
wire n_1751;
wire n_1752;
wire n_1753;
wire n_1893;
wire n_1880;
wire n_1756;
wire n_1882;
wire n_1758;
wire n_1759;
wire n_1877;
wire n_1878;
wire n_1764;
wire n_1765;
wire n_1766;
wire n_1767;
wire n_1768;
wire n_1769;
wire n_1770;
wire n_1771;
wire n_1772;
wire n_1773;
wire n_1774;
wire n_1775;
wire n_1776;
wire n_1777;
wire n_1778;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1891;
wire n_1889;
wire n_1890;
wire n_1798;
wire n_1718;
wire n_1799;
wire n_1800;
wire n_1801;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1719;
wire n_1816;
wire n_1817;
wire n_1818;
wire n_1819;
wire n_1820;
wire n_1835;
wire n_1535;
wire n_1836;
wire n_1806;
wire n_1805;
wire n_1854;
wire n_1855;
wire n_1856;
wire n_1857;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1861;
wire n_1862;
wire n_1863;
wire n_1864;
wire n_1865;
wire n_1866;
wire n_1867;
wire n_1898;
wire n_1899;
wire n_1793;
wire n_1900;
wire n_1901;
wire n_1902;
wire n_1903;
wire n_1904;
wire n_1935;
wire n_1931;
wire n_1919;
wire n_1914;
wire n_1910;
wire n_1937;
wire n_1938;
wire n_1939;
wire n_1940;
wire n_1892;
wire n_1942;
wire n_1943;
wire n_1944;
wire n_1945;
wire n_1946;
wire n_1947;
wire n_1948;
wire n_1949;
wire n_1950;
wire n_2064;
wire n_2066;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1812;
wire n_1794;
wire n_1972;
wire n_1973;
wire n_1895;
wire n_1930;
wire n_1983;
wire n_2119;
wire n_1964;
wire n_1989;
wire n_2131;
wire n_2130;
wire n_1993;
wire n_1994;
wire n_1995;
wire n_1929;
wire n_1996;
wire n_1997;
wire n_1998;
wire n_1999;
wire n_2000;
wire n_2001;
wire n_2002;
wire n_1840;
wire n_2132;
wire n_2004;
wire n_2005;
wire n_2006;
wire n_1821;
wire n_2007;
wire n_1823;
wire n_1814;
wire n_1815;
wire n_2008;
wire n_2009;
wire n_1912;
wire n_558;
wire n_1848;
wire n_256;
wire n_2010;
wire n_1928;
wire n_1926;
wire n_1925;
wire n_2011;
wire n_2012;
wire n_1837;
wire n_1838;
wire n_1841;
wire n_2013;
wire n_2014;
wire n_2015;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_2020;
wire n_2021;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2060;
wire n_2053;
wire n_2052;
wire n_2027;
wire n_1894;
wire n_2028;
wire n_2029;
wire n_2030;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2125;
wire n_2118;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2045;
wire n_2046;
wire n_2047;
wire n_2048;
wire n_2049;
wire n_2050;
wire n_2051;
wire n_2068;
wire n_2071;
wire n_2089;
wire n_2090;
wire n_2091;
wire n_2092;
wire n_2093;
wire n_2094;
wire n_2095;
wire n_2096;
wire n_2097;
wire n_2098;
wire n_2099;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2212;
wire n_2211;
wire n_2112;
wire n_2113;
wire n_2217;
wire n_2218;
wire n_2120;
wire n_2121;
wire n_2081;
wire n_2080;
wire n_2138;
wire n_2139;
wire n_2140;
wire n_2141;
wire n_2144;
wire n_2086;
wire n_2111;
wire n_2155;
wire n_1976;
wire n_1981;
wire n_1962;
wire n_1975;
wire n_2156;
wire n_2157;
wire n_1984;
wire n_2158;
wire n_1991;
wire n_2038;
wire n_1990;
wire n_2159;
wire n_2160;
wire n_2161;
wire n_2073;
wire n_2162;
wire n_2163;
wire n_2164;
wire n_2165;
wire n_2166;
wire n_2167;
wire n_2168;
wire n_2169;
wire n_2170;
wire n_2171;
wire n_2194;
wire n_2179;
wire n_2189;
wire n_2190;
wire n_2191;
wire n_2110;
wire n_2192;
wire n_2107;
wire n_2087;
wire n_2109;
wire n_2193;
wire n_2246;
wire n_2248;
wire n_2197;
wire n_2198;
wire n_2253;
wire n_2256;
wire n_2203;
wire n_2204;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2208;
wire n_2085;
wire n_2076;
wire n_2219;
wire n_2220;
wire n_2221;
wire n_2222;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2216;
wire n_2230;
wire n_2196;
wire n_2231;
wire n_2195;
wire n_2210;
wire n_2232;
wire n_2260;
wire n_2261;
wire n_2237;
wire n_2238;
wire n_2239;
wire n_2240;
wire n_2241;
wire n_2496;
wire n_2495;
wire n_2247;
wire n_2501;
wire n_2500;
wire n_2254;
wire n_2255;
wire n_2486;
wire n_2485;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2265;
wire n_2074;
wire n_2282;
wire n_2283;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2288;
wire n_2289;
wire n_2290;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2294;
wire n_2146;
wire n_2135;
wire n_2148;
wire n_2147;
wire n_2295;
wire n_2296;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_2178;
wire n_2300;
wire n_2133;
wire n_2075;
wire n_2134;
wire n_2301;
wire n_2275;
wire n_2313;
wire n_2281;
wire n_2315;
wire n_2280;
wire n_2321;
wire n_2490;
wire n_2484;
wire n_2328;
wire n_2481;
wire n_2480;
wire n_2334;
wire n_2457;
wire n_2458;
wire n_2506;
wire n_2342;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2346;
wire n_2347;
wire n_2348;
wire n_2349;
wire n_2350;
wire n_2351;
wire n_2352;
wire n_2455;
wire n_2454;
wire n_2358;
wire n_2302;
wire n_2359;
wire n_2467;
wire n_2466;
wire n_2365;
wire n_2366;
wire n_2367;
wire n_2368;
wire n_2369;
wire n_2336;
wire n_2335;
wire n_2375;
wire n_2326;
wire n_2325;
wire n_2379;
wire n_2380;
wire n_2341;
wire n_2340;
wire n_2385;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2391;
wire n_2392;
wire n_2393;
wire n_2394;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_2303;
wire n_2401;
wire n_2402;
wire n_2450;
wire n_2449;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2462;
wire n_2461;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire n_2439;
wire n_2440;
wire n_2441;
wire n_2460;
wire n_2445;
wire n_2452;
wire n_2417;
wire n_2407;
wire n_2470;
wire n_2471;
wire n_2472;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2444;
wire n_2382;
wire n_2509;
wire n_2510;
wire n_2511;
wire n_2512;
wire n_2405;
wire n_2383;
wire n_2513;
wire n_2423;
wire n_2514;
wire n_2428;
wire n_2427;
wire n_2515;
wire n_2357;
wire n_2522;
wire n_2587;
wire n_2370;
wire n_2527;
wire n_2528;
wire n_2526;
wire n_2521;
wire n_2534;
wire n_2535;
wire n_2536;
wire n_2537;
wire n_2400;
wire n_2384;
wire n_2403;
wire n_2404;
wire n_2538;
wire n_2539;
wire n_2406;
wire n_2540;
wire n_2420;
wire n_2421;
wire n_2304;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_2548;
wire n_2549;
wire n_2550;
wire n_2551;
wire n_2552;
wire n_2553;
wire n_2590;
wire n_2584;
wire n_2572;
wire n_2371;
wire n_2360;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2578;
wire n_2579;
wire n_2592;
wire n_2583;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2580;
wire n_0;
wire n_2582;
wire n_2581;
wire n_1;
wire n_2;
wire n_4;
wire n_5;
wire n_2520;
wire n_2562;
wire n_2517;
wire n_2519;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_2569;
wire n_12;
wire n_2570;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_22;
wire n_21;
wire n_27;
wire n_24;
wire n_23;
wire n_26;
wire n_113;
wire n_139;
wire n_140;
wire n_142;
wire n_146;
wire n_147;
wire n_148;
wire n_151;
wire n_166;
wire n_167;
wire n_175;
wire n_176;
wire n_181;
wire n_182;
wire n_187;
wire n_188;
wire n_204;
wire n_205;
wire n_206;
wire n_209;
wire n_226;
wire n_227;
wire n_228;
wire n_230;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_264;
wire n_265;
wire n_266;
wire n_272;
wire n_279;
wire n_277;
wire n_278;
wire n_282;
wire n_280;
wire n_313;
wire n_339;
wire n_308;
wire n_311;
wire n_319;
wire n_314;
wire n_323;
wire n_320;
wire n_326;
wire n_324;
wire n_330;
wire n_325;
wire n_328;
wire n_327;
wire n_335;
wire n_333;
wire n_332;
wire n_334;
wire n_338;
wire n_357;
wire n_356;
wire n_368;
wire n_372;
wire n_379;
wire n_377;
wire n_378;
wire n_396;
wire n_384;
wire n_382;
wire n_398;
wire n_395;
wire n_394;
wire n_400;
wire n_399;
wire n_419;
wire n_418;
wire n_420;
wire n_441;
wire n_438;
wire n_444;
wire n_442;
wire n_457;
wire n_453;
wire n_496;
wire n_488;
wire n_487;
wire n_468;
wire n_467;
wire n_557;
wire n_469;
wire n_494;
wire n_501;
wire n_498;
wire n_533;
wire n_532;
wire n_530;
wire n_515;
wire n_521;
wire n_522;
wire n_559;
wire n_531;
wire n_536;
wire n_555;
wire n_543;
wire n_535;
wire n_542;
wire n_544;
wire n_561;
wire n_562;
wire n_564;
wire n_567;
wire n_570;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_577;
wire n_583;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_608;
wire n_609;
wire n_612;
wire n_613;
wire n_616;
wire n_640;
wire n_645;
wire n_647;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_695;
wire n_696;
wire n_726;
wire n_731;
wire n_737;
wire n_762;
wire n_763;
wire n_769;
wire n_770;
wire n_771;
wire n_774;
wire n_775;
wire n_776;
wire n_778;
wire n_779;
wire n_780;
wire n_784;
wire n_817;
wire n_829;
wire n_830;
wire n_836;
wire n_835;
wire n_838;
wire n_837;
wire n_839;
wire n_842;
wire n_845;
wire n_853;
wire n_850;
wire n_852;
wire n_851;
wire n_856;
wire n_857;
wire n_885;
wire n_886;
wire n_897;
wire n_898;
wire n_943;
wire n_941;
wire n_927;
wire n_925;
wire n_910;
wire n_911;
wire n_929;
wire n_926;
wire n_1003;
wire n_1002;
wire n_938;
wire n_988;
wire n_942;
wire n_985;
wire n_987;
wire n_986;
wire n_1001;
wire n_1000;
wire n_946;
wire n_953;
wire n_952;
wire n_951;
wire n_1028;
wire n_993;
wire n_954;
wire n_984;
wire n_992;
wire n_998;
wire n_991;
wire n_996;
wire n_1027;
wire n_1004;
wire n_1006;
wire n_1005;
wire n_1007;
wire n_1015;
wire n_1009;
wire n_1024;
wire n_1018;
wire n_1014;
wire n_1016;
wire n_1023;
wire n_1026;
wire n_1025;
wire n_1034;
wire n_1033;
wire n_1049;
wire n_1055;
wire n_1054;
wire n_1057;
wire n_1065;
wire n_1064;
wire n_1058;
wire n_1059;
wire n_1102;
wire n_1101;
wire n_1100;
wire n_1098;
wire n_1095;
wire n_1111;
wire n_1104;
wire n_1099;
wire n_1110;
wire n_1119;
wire n_1118;
wire n_1112;
wire n_1129;
wire n_1143;
wire n_1121;
wire n_1122;
wire n_1197;
wire n_1146;
wire n_1153;
wire n_1147;
wire n_1152;
wire n_1151;
wire n_1190;
wire n_1154;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1164;
wire n_1194;
wire n_1193;
wire n_1212;
wire n_1198;
wire n_1205;
wire n_1203;
wire n_1204;
wire n_1222;
wire n_1213;
wire n_1228;
wire n_1227;
wire n_1230;
wire n_1262;
wire n_1261;
wire n_1294;
wire n_1293;
wire n_1266;
wire n_1290;
wire n_1291;
wire n_1299;
wire n_1303;
wire n_1297;
wire n_1298;
wire n_1302;
wire n_1305;
wire n_1320;
wire n_1322;
wire n_1324;
wire n_1325;
wire n_1328;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1343;
wire n_1345;
wire n_1346;
wire n_1348;
wire n_1349;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1363;
wire n_1364;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1373;
wire n_1374;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1414;
wire n_1415;
wire n_1419;
wire n_1421;
wire n_1422;
wire n_1424;
wire n_1425;
wire n_1447;
wire n_1453;
wire n_1452;
wire n_1455;
wire n_1454;
wire n_1477;
wire n_1476;
wire n_1533;
wire n_1459;
wire n_1456;
wire n_1460;
wire n_1480;
wire n_1483;
wire n_1531;
wire n_1506;
wire n_1507;
wire n_1524;
wire n_1523;
wire n_1529;
wire n_1527;
wire n_1528;
wire n_1574;
wire n_1553;
wire n_1563;
wire n_1554;
wire n_1557;
wire n_1555;
wire n_1560;
wire n_1558;
wire n_1562;
wire n_1561;
wire n_1559;
wire n_1567;
wire n_1566;
wire n_1569;
wire n_1568;
wire n_1610;
wire n_1609;
wire n_1608;
wire n_1575;
wire n_1586;
wire n_1580;
wire n_1579;
wire n_1576;
wire n_1577;
wire n_1590;
wire n_1588;
wire n_1607;
wire n_1589;
wire n_1603;
wire n_1606;
wire n_1605;
wire n_1649;
wire n_1613;
wire n_1622;
wire n_1621;
wire n_1614;
wire n_1617;
wire n_1620;
wire n_1624;
wire n_1623;
wire n_1629;
wire n_1647;
wire n_1634;
wire n_1628;
wire n_1630;
wire n_1640;
wire n_1650;
wire n_1652;
wire n_1653;
wire n_1654;
wire n_1659;
wire n_1660;
wire n_1661;
wire n_1698;
wire n_1699;
wire n_1700;
wire n_1701;
wire n_1702;
wire n_1703;
wire n_1704;
wire n_1705;
wire n_1706;
wire n_1707;
wire n_1708;
wire n_1709;
wire n_1712;
wire n_1713;
wire n_1714;
wire n_1715;
wire n_1716;
wire n_1757;
wire n_1720;
wire n_1728;
wire n_1721;
wire n_1723;
wire n_1722;
wire n_1725;
wire n_1724;
wire n_1783;
wire n_1726;
wire n_1737;
wire n_1736;
wire n_1732;
wire n_1790;
wire n_1733;
wire n_1740;
wire n_1744;
wire n_1743;
wire n_1755;
wire n_1754;
wire n_1785;
wire n_1761;
wire n_1763;
wire n_1782;
wire n_1789;
wire n_1796;
wire n_1795;
wire n_1811;
wire n_1797;
wire n_1807;
wire n_1845;
wire n_1844;
wire n_1810;
wire n_1808;
wire n_1851;
wire n_1809;
wire n_1869;
wire n_1868;
wire n_1832;
wire n_1813;
wire n_1822;
wire n_1875;
wire n_1830;
wire n_1829;
wire n_1828;
wire n_1824;
wire n_1827;
wire n_1826;
wire n_1831;
wire n_1842;
wire n_1833;
wire n_1834;
wire n_1839;
wire n_1849;
wire n_1843;
wire n_1846;
wire n_1847;
wire n_1853;
wire n_1850;
wire n_1852;
wire n_1870;
wire n_1872;
wire n_1871;
wire n_1873;
wire n_1874;
wire n_1876;
wire n_1879;
wire n_1883;
wire n_1884;
wire n_1885;
wire n_1886;
wire n_1887;
wire n_1888;
wire n_1896;
wire n_1905;
wire n_1897;
wire n_1907;
wire n_1906;
wire n_1915;
wire n_1954;
wire n_1951;
wire n_1941;
wire n_1909;
wire n_1908;
wire n_1923;
wire n_1918;
wire n_1911;
wire n_1913;
wire n_1917;
wire n_1916;
wire n_1921;
wire n_1920;
wire n_1922;
wire n_1924;
wire n_1927;
wire n_1952;
wire n_1936;
wire n_1932;
wire n_1934;
wire n_1933;
wire n_1953;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1963;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1974;
wire n_1977;
wire n_1978;
wire n_1979;
wire n_1980;
wire n_1982;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1988;
wire n_1992;
wire n_2003;
wire n_2025;
wire n_2026;
wire n_2037;
wire n_2039;
wire n_2040;
wire n_2041;
wire n_2054;
wire n_2055;
wire n_2056;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_2061;
wire n_2062;
wire n_2063;
wire n_2065;
wire n_2067;
wire n_2069;
wire n_2070;
wire n_2072;
wire n_2077;
wire n_2079;
wire n_2078;
wire n_2082;
wire n_2149;
wire n_2175;
wire n_2174;
wire n_2084;
wire n_2083;
wire n_2153;
wire n_2152;
wire n_2200;
wire n_2114;
wire n_2088;
wire n_2108;
wire n_2236;
wire n_2116;
wire n_2115;
wire n_2126;
wire n_2117;
wire n_2124;
wire n_2122;
wire n_2123;
wire n_2129;
wire n_2127;
wire n_2128;
wire n_2234;
wire n_2137;
wire n_2136;
wire n_2143;
wire n_2142;
wire n_2145;
wire n_2215;
wire n_2184;
wire n_2183;
wire n_2182;
wire n_2150;
wire n_2173;
wire n_2151;
wire n_2177;
wire n_2154;
wire n_2172;
wire n_2176;
wire n_2181;
wire n_2180;
wire n_2186;
wire n_2185;
wire n_2188;
wire n_2209;
wire n_2187;
wire n_2199;
wire n_2201;
wire n_2202;
wire n_2213;
wire n_2214;
wire n_2235;
wire n_2233;
wire n_2242;
wire n_2244;
wire n_2245;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2266;
wire n_2267;
wire n_2268;
wire n_2269;
wire n_2270;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2276;
wire n_2277;
wire n_2278;
wire n_2279;
wire n_2305;
wire n_2307;
wire n_2322;
wire n_2306;
wire n_2310;
wire n_2308;
wire n_2309;
wire n_2355;
wire n_2320;
wire n_2319;
wire n_2318;
wire n_2316;
wire n_2312;
wire n_2311;
wire n_2314;
wire n_2327;
wire n_2317;
wire n_2331;
wire n_2330;
wire n_2323;
wire n_2324;
wire n_2329;
wire n_2333;
wire n_2332;
wire n_2339;
wire n_2356;
wire n_2337;
wire n_2338;
wire n_2353;
wire n_2354;
wire n_2363;
wire n_2361;
wire n_2364;
wire n_2362;
wire n_2372;
wire n_2377;
wire n_2374;
wire n_2373;
wire n_2376;
wire n_2381;
wire n_2378;
wire n_2430;
wire n_2410;
wire n_2408;
wire n_2419;
wire n_2418;
wire n_2409;
wire n_2413;
wire n_2443;
wire n_2411;
wire n_2412;
wire n_2425;
wire n_2424;
wire n_2433;
wire n_2432;
wire n_2422;
wire n_2431;
wire n_2429;
wire n_2426;
wire n_2442;
wire n_2446;
wire n_2448;
wire n_2447;
wire n_2453;
wire n_2451;
wire n_2456;
wire n_2505;
wire n_2459;
wire n_2507;
wire n_2504;
wire n_2463;
wire n_2465;
wire n_2464;
wire n_2468;
wire n_2479;
wire n_2469;
wire n_2494;
wire n_2493;
wire n_2491;
wire n_2483;
wire n_2482;
wire n_2516;
wire n_2508;
wire n_2487;
wire n_2489;
wire n_2488;
wire n_2492;
wire n_2502;
wire n_2499;
wire n_2497;
wire n_2498;
wire n_2503;
wire n_2518;
wire n_2523;
wire n_2524;
wire n_2525;
wire n_2529;
wire n_2530;
wire n_2531;
wire n_2532;
wire n_2533;
wire n_2541;
wire n_2554;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2561;
wire n_2563;
wire n_2564;
wire n_2565;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2571;
wire n_2593;
wire n_2586;
wire n_2585;
wire n_2588;
wire n_2589;
wire n_2591;
wire n_2600;
wire n_2599;
wire n_2598;


INV_X1 i_2629 (.ZN (n_2600), .A (n_2533));
XNOR2_X1 i_2628 (.ZN (n_2599), .A (n_2559), .B (n_2523));
XOR2_X1 i_2627 (.Z (n_2598), .A (n_2571), .B (n_2518));
NAND2_X1 i_2626 (.ZN (n_2593), .A1 (n_2599), .A2 (n_2598));
OAI21_X1 i_2625 (.ZN (n_2592), .A (n_2593), .B1 (n_2599), .B2 (n_2598));
NOR2_X1 i_2624 (.ZN (n_2591), .A1 (n_2531), .A2 (n_2600));
XNOR2_X1 i_2623 (.ZN (n_2590), .A (n_2532), .B (n_2591));
NOR2_X1 i_2613 (.ZN (n_2589), .A1 (n_2361), .A2 (n_2541));
AOI22_X1 i_2612 (.ZN (n_2588), .A1 (A[20]), .A2 (B[21]), .B1 (A[19]), .B2 (B[22]));
NOR2_X1 i_2611 (.ZN (n_2587), .A1 (n_2589), .A2 (n_2588));
OAI22_X1 i_2610 (.ZN (n_2586), .A1 (n_2361), .A2 (n_2541), .B1 (n_2370), .B2 (n_2588));
XOR2_X1 i_2609 (.Z (n_2585), .A (n_2555), .B (n_2556));
XOR2_X1 i_2608 (.Z (n_2584), .A (n_2586), .B (n_2585));
AOI22_X1 i_2607 (.ZN (n_2583), .A1 (n_2586), .A2 (n_2585), .B1 (n_2590), .B2 (n_2584));
OAI21_X1 i_2606 (.ZN (n_2582), .A (n_2593), .B1 (n_2592), .B2 (n_2583));
XNOR2_X1 i_2605 (.ZN (n_2581), .A (n_2561), .B (n_2568));
NAND2_X1 i_2604 (.ZN (n_2580), .A1 (n_2582), .A2 (n_2581));
NOR2_X1 i_2603 (.ZN (n_2571), .A1 (n_2566), .A2 (n_2564));
INV_X1 i_2602 (.ZN (n_2570), .A (n_2569));
AOI22_X1 i_2601 (.ZN (n_2569), .A1 (n_2561), .A2 (n_2568), .B1 (n_2563), .B2 (n_2567));
XOR2_X1 i_2600 (.Z (n_2568), .A (n_2563), .B (n_2567));
OAI21_X1 i_2599 (.ZN (n_2567), .A (n_2565), .B1 (n_2566), .B2 (n_2518));
NOR2_X1 i_2598 (.ZN (n_2566), .A1 (n_2554), .A2 (n_2517));
INV_X1 i_2597 (.ZN (n_2565), .A (n_2564));
AOI22_X1 i_2596 (.ZN (n_2564), .A1 (A[21]), .A2 (B[22]), .B1 (B[21]), .B2 (A[22]));
XNOR2_X1 i_2590 (.ZN (n_2563), .A (n_2520), .B (n_2562));
NAND2_X1 i_2586 (.ZN (n_2562), .A1 (B[21]), .A2 (A[23]));
AOI22_X1 i_2585 (.ZN (n_2561), .A1 (n_2559), .A2 (n_2560), .B1 (n_2557), .B2 (n_2558));
INV_X1 i_2584 (.ZN (n_2560), .A (n_2523));
XOR2_X1 i_2583 (.Z (n_2559), .A (n_2557), .B (n_2558));
OAI22_X1 i_2582 (.ZN (n_2558), .A1 (n_2555), .A2 (n_2556), .B1 (n_2554), .B2 (n_2541));
AOI21_X1 i_2581 (.ZN (n_2557), .A (n_2531), .B1 (n_2532), .B2 (n_2533));
NAND2_X1 i_2580 (.ZN (n_2556), .A1 (B[23]), .A2 (A[19]));
XNOR2_X1 i_2579 (.ZN (n_2555), .A (n_2554), .B (n_2541));
NAND2_X1 i_2578 (.ZN (n_2554), .A1 (B[21]), .A2 (A[21]));
NAND2_X1 i_2577 (.ZN (n_2541), .A1 (B[22]), .A2 (A[20]));
NAND3_X1 i_2576 (.ZN (n_2533), .A1 (n_2530), .A2 (B[19]), .A3 (A[23]));
NAND2_X1 i_2575 (.ZN (n_2532), .A1 (B[20]), .A2 (A[22]));
AOI21_X1 i_2574 (.ZN (n_2531), .A (n_2530), .B1 (B[19]), .B2 (A[23]));
NAND2_X1 i_2573 (.ZN (n_2530), .A1 (n_2528), .A2 (n_2529));
INV_X1 i_2572 (.ZN (n_2529), .A (n_2524));
NAND2_X1 i_2571 (.ZN (n_2528), .A1 (n_2526), .A2 (n_2521));
NOR2_X1 i_2570 (.ZN (n_2526), .A1 (n_2524), .A2 (n_2525));
AOI22_X1 i_2569 (.ZN (n_2525), .A1 (A[21]), .A2 (B[20]), .B1 (B[18]), .B2 (A[23]));
NOR2_X1 i_2568 (.ZN (n_2524), .A1 (n_2523), .A2 (n_2381));
NAND2_X1 i_2567 (.ZN (n_2523), .A1 (B[20]), .A2 (A[23]));
INV_X1 i_2566 (.ZN (n_2521), .A (n_2378));
XNOR2_X1 i_2565 (.ZN (n_2520), .A (n_2517), .B (n_2519));
NAND2_X1 i_2564 (.ZN (n_2519), .A1 (A[21]), .A2 (B[23]));
NOR2_X1 i_2563 (.ZN (n_2518), .A1 (n_1322), .A2 (n_1533));
NAND2_X1 i_2562 (.ZN (n_2517), .A1 (A[22]), .A2 (B[22]));
INV_X1 i_2561 (.ZN (n_2516), .A (A[14]));
INV_X1 i_2560 (.ZN (n_2508), .A (B[21]));
INV_X1 i_2559 (.ZN (n_2507), .A (n_2340));
INV_X1 i_2558 (.ZN (n_2506), .A (n_2356));
NAND2_X1 i_2557 (.ZN (n_2505), .A1 (A[16]), .A2 (B[19]));
INV_X1 i_2556 (.ZN (n_2504), .A (n_2505));
NOR2_X1 i_2555 (.ZN (n_2503), .A1 (n_558), .A2 (n_856));
NAND2_X1 i_2554 (.ZN (n_2502), .A1 (n_2504), .A2 (n_2503));
OAI21_X1 i_2553 (.ZN (n_2501), .A (n_2502), .B1 (n_2504), .B2 (n_2503));
NAND2_X1 i_2552 (.ZN (n_2500), .A1 (A[17]), .A2 (B[18]));
OR2_X1 i_2550 (.ZN (n_2499), .A1 (n_2249), .A2 (n_2266));
AOI22_X1 i_2549 (.ZN (n_2498), .A1 (A[19]), .A2 (B[16]), .B1 (A[20]), .B2 (B[15]));
INV_X1 i_2548 (.ZN (n_2497), .A (n_2498));
NAND2_X1 i_2547 (.ZN (n_2496), .A1 (n_2499), .A2 (n_2497));
NAND2_X1 i_2546 (.ZN (n_2495), .A1 (A[18]), .A2 (B[17]));
OAI21_X1 i_2545 (.ZN (n_2494), .A (n_2499), .B1 (n_2496), .B2 (n_2495));
OAI21_X1 i_2544 (.ZN (n_2493), .A (n_2502), .B1 (n_2501), .B2 (n_2500));
NAND2_X1 i_2543 (.ZN (n_2492), .A1 (n_2494), .A2 (n_2493));
INV_X1 i_2542 (.ZN (n_2491), .A (n_2492));
OAI21_X1 i_2541 (.ZN (n_2490), .A (n_2492), .B1 (n_2494), .B2 (n_2493));
NOR2_X1 i_2540 (.ZN (n_2489), .A1 (n_2516), .A2 (n_2508));
NOR2_X1 i_2539 (.ZN (n_2488), .A1 (n_256), .A2 (n_1368));
NAND2_X1 i_2538 (.ZN (n_2487), .A1 (n_2489), .A2 (n_2488));
OAI21_X1 i_2537 (.ZN (n_2486), .A (n_2487), .B1 (n_2489), .B2 (n_2488));
NAND2_X1 i_2536 (.ZN (n_2485), .A1 (A[12]), .A2 (B[23]));
OAI21_X1 i_2535 (.ZN (n_2484), .A (n_2487), .B1 (n_2486), .B2 (n_2485));
NOR3_X1 i_2534 (.ZN (n_2483), .A1 (n_2516), .A2 (n_2508), .A3 (n_2329));
AOI22_X1 i_2533 (.ZN (n_2482), .A1 (A[14]), .A2 (B[22]), .B1 (A[15]), .B2 (B[21]));
NOR2_X1 i_2532 (.ZN (n_2481), .A1 (n_2483), .A2 (n_2482));
NOR2_X1 i_2531 (.ZN (n_2480), .A1 (n_256), .A2 (n_1533));
AOI21_X1 i_2530 (.ZN (n_2479), .A (n_2483), .B1 (n_2481), .B2 (n_2480));
OAI22_X1 i_2529 (.ZN (n_2469), .A1 (n_2494), .A2 (n_2493), .B1 (n_2491), .B2 (n_2484));
NOR2_X1 i_2528 (.ZN (n_2468), .A1 (n_2479), .A2 (n_2469));
AOI21_X1 i_2527 (.ZN (n_2467), .A (n_2468), .B1 (n_2479), .B2 (n_2469));
OAI22_X1 i_2526 (.ZN (n_2466), .A1 (n_2279), .A2 (n_2278), .B1 (n_2276), .B2 (n_2277));
AOI21_X1 i_2525 (.ZN (n_2465), .A (n_2468), .B1 (n_2467), .B2 (n_2466));
XNOR2_X1 i_2524 (.ZN (n_2464), .A (n_2312), .B (n_2311));
NOR2_X1 i_2523 (.ZN (n_2463), .A1 (n_2465), .A2 (n_2464));
AOI21_X1 i_2522 (.ZN (n_2462), .A (n_2463), .B1 (n_2465), .B2 (n_2464));
XNOR2_X1 i_2521 (.ZN (n_2461), .A (n_2330), .B (n_2324));
AOI21_X1 i_2520 (.ZN (n_2460), .A (n_2463), .B1 (n_2462), .B2 (n_2461));
AOI22_X1 i_2519 (.ZN (n_2459), .A1 (A[17]), .A2 (B[19]), .B1 (A[16]), .B2 (B[20]));
AOI21_X1 i_2518 (.ZN (n_2458), .A (n_2459), .B1 (n_2507), .B2 (n_2504));
NAND2_X1 i_2517 (.ZN (n_2457), .A1 (n_2506), .A2 (n_2458));
OAI21_X1 i_2516 (.ZN (n_2456), .A (n_2457), .B1 (n_2340), .B2 (n_2505));
XOR2_X1 i_2514 (.Z (n_2455), .A (n_2145), .B (n_2456));
OAI21_X1 i_2513 (.ZN (n_2454), .A (n_2269), .B1 (n_2271), .B2 (n_2272));
AOI22_X1 i_2512 (.ZN (n_2453), .A1 (n_2145), .A2 (n_2456), .B1 (n_2455), .B2 (n_2454));
XNOR2_X1 i_2511 (.ZN (n_2451), .A (n_2319), .B (n_2318));
XOR2_X1 i_2510 (.Z (n_2450), .A (n_2453), .B (n_2451));
XOR2_X1 i_2509 (.Z (n_2449), .A (n_2411), .B (n_2339));
AOI22_X1 i_2508 (.ZN (n_2448), .A1 (n_2453), .A2 (n_2451), .B1 (n_2450), .B2 (n_2449));
XOR2_X1 i_2507 (.Z (n_2447), .A (n_2322), .B (n_2306));
NOR2_X1 i_2506 (.ZN (n_2446), .A1 (n_2448), .A2 (n_2447));
AOI21_X1 i_2505 (.ZN (n_2445), .A (n_2446), .B1 (n_2448), .B2 (n_2447));
AOI21_X1 i_2504 (.ZN (n_2444), .A (n_2446), .B1 (n_2460), .B2 (n_2445));
INV_X1 i_2503 (.ZN (n_2443), .A (n_2339));
NAND2_X1 i_2502 (.ZN (n_2442), .A1 (A[18]), .A2 (B[21]));
XNOR2_X1 i_2501 (.ZN (n_2433), .A (n_2317), .B (n_2442));
NAND2_X1 i_2500 (.ZN (n_2432), .A1 (A[16]), .A2 (B[23]));
OAI22_X1 i_2499 (.ZN (n_2431), .A1 (n_2317), .A2 (n_2442), .B1 (n_2433), .B2 (n_2432));
NAND2_X1 i_2498 (.ZN (n_2430), .A1 (A[23]), .A2 (B[17]));
INV_X1 i_2497 (.ZN (n_2429), .A (n_2430));
NOR2_X1 i_2496 (.ZN (n_2428), .A1 (n_2431), .A2 (n_2429));
NAND2_X1 i_2495 (.ZN (n_2427), .A1 (n_2431), .A2 (n_2429));
NAND2_X1 i_2494 (.ZN (n_2426), .A1 (A[20]), .A2 (B[19]));
XNOR2_X1 i_2493 (.ZN (n_2425), .A (n_2381), .B (n_2426));
NAND2_X1 i_2492 (.ZN (n_2424), .A1 (A[19]), .A2 (B[20]));
OAI22_X1 i_2491 (.ZN (n_2423), .A1 (n_2381), .A2 (n_2426), .B1 (n_2425), .B2 (n_2424));
AOI21_X1 i_2490 (.ZN (n_2422), .A (n_2428), .B1 (n_2431), .B2 (n_2429));
XOR2_X1 i_2489 (.Z (n_2421), .A (n_2423), .B (n_2422));
XNOR2_X1 i_2488 (.ZN (n_2420), .A (n_2305), .B (n_2421));
XOR2_X1 i_2487 (.Z (n_2419), .A (n_2433), .B (n_2432));
XOR2_X1 i_2486 (.Z (n_2418), .A (n_2425), .B (n_2424));
XOR2_X1 i_2485 (.Z (n_2417), .A (n_2419), .B (n_2418));
NOR2_X1 i_2484 (.ZN (n_2413), .A1 (n_2267), .A2 (n_2430));
AOI22_X1 i_2483 (.ZN (n_2412), .A1 (A[23]), .A2 (B[15]), .B1 (A[21]), .B2 (B[17]));
NOR2_X1 i_2482 (.ZN (n_2411), .A1 (n_2413), .A2 (n_2412));
AOI21_X1 i_2481 (.ZN (n_2410), .A (n_2413), .B1 (n_2443), .B2 (n_2411));
OAI22_X1 i_2480 (.ZN (n_2409), .A1 (n_1232), .A2 (n_1881), .B1 (n_592), .B2 (n_1792));
OAI21_X1 i_2476 (.ZN (n_2408), .A (n_2409), .B1 (n_2339), .B2 (n_2430));
XOR2_X1 i_2475 (.Z (n_2407), .A (n_2410), .B (n_2408));
AOI22_X1 i_2474 (.ZN (n_2406), .A1 (n_2419), .A2 (n_2418), .B1 (n_2417), .B2 (n_2407));
XNOR2_X1 i_2473 (.ZN (n_2405), .A (n_2420), .B (n_2406));
XOR2_X1 i_2472 (.Z (n_2404), .A (n_2374), .B (n_2373));
OAI22_X1 i_2471 (.ZN (n_2403), .A1 (n_2339), .A2 (n_2430), .B1 (n_2410), .B2 (n_2408));
XOR2_X1 i_2470 (.Z (n_2400), .A (n_2404), .B (n_2403));
XNOR2_X1 i_2469 (.ZN (n_2384), .A (n_2362), .B (n_2361));
XOR2_X1 i_2468 (.Z (n_2383), .A (n_2400), .B (n_2384));
XOR2_X1 i_2467 (.Z (n_2382), .A (n_2405), .B (n_2383));
NAND2_X1 i_2466 (.ZN (n_2381), .A1 (B[18]), .A2 (A[21]));
NAND2_X1 i_2465 (.ZN (n_2378), .A1 (B[19]), .A2 (A[22]));
NOR2_X1 i_2464 (.ZN (n_2377), .A1 (n_2381), .A2 (n_2378));
AOI22_X1 i_2463 (.ZN (n_2376), .A1 (B[19]), .A2 (A[21]), .B1 (B[18]), .B2 (A[22]));
NOR2_X1 i_2462 (.ZN (n_2374), .A1 (n_2377), .A2 (n_2376));
NOR2_X1 i_2461 (.ZN (n_2373), .A1 (n_1322), .A2 (n_856));
AOI21_X1 i_2460 (.ZN (n_2372), .A (n_2377), .B1 (n_2374), .B2 (n_2373));
INV_X1 i_2459 (.ZN (n_2371), .A (n_2372));
NAND2_X1 i_2458 (.ZN (n_2370), .A1 (B[23]), .A2 (A[18]));
NOR2_X1 i_2457 (.ZN (n_2364), .A1 (n_2317), .A2 (n_2370));
AOI22_X1 i_2456 (.ZN (n_2363), .A1 (B[23]), .A2 (A[17]), .B1 (B[22]), .B2 (A[18]));
NOR2_X1 i_2455 (.ZN (n_2362), .A1 (n_2364), .A2 (n_2363));
NAND2_X1 i_2454 (.ZN (n_2361), .A1 (B[21]), .A2 (A[19]));
OAI22_X1 i_2453 (.ZN (n_2360), .A1 (n_2317), .A2 (n_2370), .B1 (n_2363), .B2 (n_2361));
XOR2_X1 i_2452 (.Z (n_2357), .A (n_2371), .B (n_2360));
NAND2_X1 i_2451 (.ZN (n_2356), .A1 (A[18]), .A2 (B[18]));
NAND2_X1 i_2450 (.ZN (n_2355), .A1 (A[19]), .A2 (B[19]));
AOI22_X1 i_2449 (.ZN (n_2354), .A1 (A[18]), .A2 (B[19]), .B1 (A[19]), .B2 (B[18]));
INV_X1 i_2448 (.ZN (n_2353), .A (n_2354));
OAI21_X1 i_2447 (.ZN (n_2341), .A (n_2353), .B1 (n_2356), .B2 (n_2355));
NAND2_X1 i_2446 (.ZN (n_2340), .A1 (A[17]), .A2 (B[20]));
NAND2_X1 i_2445 (.ZN (n_2339), .A1 (A[22]), .A2 (B[16]));
AOI22_X1 i_2444 (.ZN (n_2338), .A1 (A[22]), .A2 (B[15]), .B1 (A[21]), .B2 (B[16]));
INV_X1 i_2443 (.ZN (n_2337), .A (n_2338));
OAI21_X1 i_2442 (.ZN (n_2336), .A (n_2337), .B1 (n_2267), .B2 (n_2339));
NAND2_X1 i_2441 (.ZN (n_2335), .A1 (A[20]), .A2 (B[17]));
OAI22_X1 i_2440 (.ZN (n_2333), .A1 (n_2356), .A2 (n_2355), .B1 (n_2341), .B2 (n_2340));
OAI22_X1 i_2439 (.ZN (n_2332), .A1 (n_2267), .A2 (n_2339), .B1 (n_2336), .B2 (n_2335));
NAND2_X1 i_2438 (.ZN (n_2331), .A1 (n_2333), .A2 (n_2332));
OAI21_X1 i_2437 (.ZN (n_2330), .A (n_2331), .B1 (n_2333), .B2 (n_2332));
NAND2_X1 i_2436 (.ZN (n_2329), .A1 (A[15]), .A2 (B[22]));
NAND2_X1 i_2435 (.ZN (n_2327), .A1 (A[16]), .A2 (B[21]));
XNOR2_X1 i_2434 (.ZN (n_2326), .A (n_2329), .B (n_2327));
NAND2_X1 i_2433 (.ZN (n_2325), .A1 (A[14]), .A2 (B[23]));
OAI22_X1 i_2432 (.ZN (n_2324), .A1 (n_2329), .A2 (n_2327), .B1 (n_2326), .B2 (n_2325));
INV_X1 i_2430 (.ZN (n_2323), .A (n_2324));
OAI21_X1 i_2429 (.ZN (n_2322), .A (n_2331), .B1 (n_2330), .B2 (n_2323));
NAND2_X1 i_2428 (.ZN (n_2320), .A1 (A[20]), .A2 (B[18]));
XNOR2_X1 i_2427 (.ZN (n_2319), .A (n_2355), .B (n_2320));
NAND2_X1 i_2426 (.ZN (n_2318), .A1 (A[18]), .A2 (B[20]));
NAND2_X1 i_2425 (.ZN (n_2317), .A1 (A[17]), .A2 (B[22]));
NOR2_X1 i_2424 (.ZN (n_2316), .A1 (n_2327), .A2 (n_2317));
AOI22_X1 i_2423 (.ZN (n_2314), .A1 (A[16]), .A2 (B[22]), .B1 (A[17]), .B2 (B[21]));
NOR2_X1 i_2422 (.ZN (n_2312), .A1 (n_2316), .A2 (n_2314));
NOR2_X1 i_2421 (.ZN (n_2311), .A1 (n_558), .A2 (n_1533));
AOI21_X1 i_2420 (.ZN (n_2310), .A (n_2316), .B1 (n_2312), .B2 (n_2311));
OAI22_X1 i_2419 (.ZN (n_2309), .A1 (n_2355), .A2 (n_2320), .B1 (n_2319), .B2 (n_2318));
INV_X1 i_2418 (.ZN (n_2308), .A (n_2309));
NOR2_X1 i_2417 (.ZN (n_2307), .A1 (n_2310), .A2 (n_2308));
AOI21_X1 i_2416 (.ZN (n_2306), .A (n_2307), .B1 (n_2310), .B2 (n_2308));
AOI21_X1 i_2415 (.ZN (n_2305), .A (n_2307), .B1 (n_2322), .B2 (n_2306));
INV_X1 i_2414 (.ZN (n_2304), .A (n_2305));
INV_X1 i_2413 (.ZN (n_2303), .A (n_2302));
AOI21_X1 i_2412 (.ZN (n_2302), .A (n_2275), .B1 (n_2281), .B2 (n_2280));
NAND2_X1 i_2411 (.ZN (n_2281), .A1 (n_2273), .A2 (n_2274));
XNOR2_X1 i_2410 (.ZN (n_2280), .A (n_2279), .B (n_2278));
XNOR2_X1 i_2409 (.ZN (n_2279), .A (n_2276), .B (n_2277));
NAND2_X1 i_2408 (.ZN (n_2278), .A1 (B[14]), .A2 (A[22]));
NAND2_X1 i_2407 (.ZN (n_2277), .A1 (B[13]), .A2 (A[23]));
AOI21_X1 i_2406 (.ZN (n_2276), .A (n_2143), .B1 (n_2137), .B2 (n_2136));
NOR2_X1 i_2405 (.ZN (n_2275), .A1 (n_2273), .A2 (n_2274));
XNOR2_X1 i_2404 (.ZN (n_2274), .A (n_2270), .B (n_2272));
OAI21_X1 i_2403 (.ZN (n_2273), .A (n_2259), .B1 (n_2260), .B2 (n_2261));
NAND2_X1 i_2402 (.ZN (n_2272), .A1 (B[17]), .A2 (A[19]));
INV_X1 i_2401 (.ZN (n_2271), .A (n_2270));
AOI21_X1 i_2400 (.ZN (n_2270), .A (n_2268), .B1 (n_2266), .B2 (n_2267));
INV_X1 i_2399 (.ZN (n_2269), .A (n_2268));
NOR2_X1 i_2398 (.ZN (n_2268), .A1 (n_2266), .A2 (n_2267));
NAND2_X1 i_2397 (.ZN (n_2267), .A1 (B[15]), .A2 (A[21]));
NAND2_X1 i_2396 (.ZN (n_2266), .A1 (B[16]), .A2 (A[20]));
AOI21_X1 i_2395 (.ZN (n_2261), .A (n_2188), .B1 (n_2186), .B2 (n_2185));
OAI21_X1 i_2394 (.ZN (n_2260), .A (n_2259), .B1 (n_2258), .B2 (n_2257));
NAND2_X1 i_2393 (.ZN (n_2259), .A1 (n_2257), .A2 (n_2258));
OAI22_X1 i_2392 (.ZN (n_2258), .A1 (n_2246), .A2 (n_2248), .B1 (n_2245), .B2 (n_2177));
OAI21_X1 i_2391 (.ZN (n_2257), .A (n_2252), .B1 (n_2253), .B2 (n_2256));
NAND2_X1 i_2390 (.ZN (n_2256), .A1 (A[17]), .A2 (B[17]));
OAI21_X1 i_2389 (.ZN (n_2253), .A (n_2252), .B1 (n_2251), .B2 (n_2250));
NAND2_X1 i_2388 (.ZN (n_2252), .A1 (n_2250), .A2 (n_2251));
INV_X1 i_2387 (.ZN (n_2251), .A (n_2249));
AND2_X1 i_2385 (.ZN (n_2250), .A1 (A[18]), .A2 (B[16]));
NAND2_X1 i_2384 (.ZN (n_2249), .A1 (B[15]), .A2 (A[19]));
NAND2_X1 i_2383 (.ZN (n_2248), .A1 (A[20]), .A2 (B[14]));
XNOR2_X1 i_2382 (.ZN (n_2246), .A (n_2245), .B (n_2177));
NAND2_X1 i_2381 (.ZN (n_2245), .A1 (B[12]), .A2 (A[22]));
INV_X1 i_2380 (.ZN (n_2244), .A (n_1966));
INV_X1 i_2379 (.ZN (n_2243), .A (B[10]));
INV_X1 i_2378 (.ZN (n_2242), .A (n_1959));
INV_X1 i_2377 (.ZN (n_2236), .A (n_1992));
OAI21_X1 i_2376 (.ZN (n_2235), .A (n_2244), .B1 (n_1967), .B2 (n_1963));
NAND2_X1 i_2375 (.ZN (n_2234), .A1 (B[12]), .A2 (A[19]));
OAI33_X1 i_2374 (.ZN (n_2233), .A1 (n_229), .A2 (n_1322), .A3 (n_2234), .B1 (n_1987)
    , .B2 (n_559), .B3 (n_1028));
XOR2_X1 i_2373 (.Z (n_2218), .A (n_2235), .B (n_2233));
AOI21_X1 i_2372 (.ZN (n_2217), .A (n_1960), .B1 (n_2242), .B2 (n_1957));
AOI22_X1 i_2371 (.ZN (n_2216), .A1 (n_2235), .A2 (n_2233), .B1 (n_2218), .B2 (n_2217));
NAND2_X1 i_2370 (.ZN (n_2215), .A1 (B[22]), .A2 (A[12]));
AOI22_X1 i_2369 (.ZN (n_2214), .A1 (B[22]), .A2 (A[11]), .B1 (B[21]), .B2 (A[12]));
INV_X1 i_2368 (.ZN (n_2213), .A (n_2214));
OAI21_X1 i_2367 (.ZN (n_2212), .A (n_2213), .B1 (n_1977), .B2 (n_2215));
NAND2_X1 i_2366 (.ZN (n_2211), .A1 (B[23]), .A2 (A[10]));
OAI22_X1 i_2365 (.ZN (n_2210), .A1 (n_1977), .A2 (n_2215), .B1 (n_2212), .B2 (n_2211));
NAND2_X1 i_2364 (.ZN (n_2209), .A1 (B[19]), .A2 (A[15]));
AOI22_X1 i_2363 (.ZN (n_2202), .A1 (B[19]), .A2 (A[14]), .B1 (B[18]), .B2 (A[15]));
INV_X1 i_2362 (.ZN (n_2201), .A (n_2202));
OAI21_X1 i_2361 (.ZN (n_2200), .A (n_2201), .B1 (n_1957), .B2 (n_2209));
OAI22_X1 i_2360 (.ZN (n_2199), .A1 (n_1957), .A2 (n_2209), .B1 (n_1958), .B2 (n_2200));
INV_X1 i_2359 (.ZN (n_2196), .A (n_2199));
XOR2_X1 i_2358 (.Z (n_2195), .A (n_2210), .B (n_2199));
XNOR2_X1 i_2357 (.ZN (n_2194), .A (n_2216), .B (n_2195));
NOR3_X1 i_2356 (.ZN (n_2188), .A1 (n_1305), .A2 (n_2209), .A3 (n_1532));
NAND2_X1 i_2355 (.ZN (n_2187), .A1 (B[18]), .A2 (A[16]));
AOI21_X1 i_2354 (.ZN (n_2186), .A (n_2188), .B1 (n_2209), .B2 (n_2187));
NOR2_X1 i_2353 (.ZN (n_2185), .A1 (n_557), .A2 (n_856));
NAND2_X1 i_2352 (.ZN (n_2184), .A1 (B[21]), .A2 (A[13]));
XNOR2_X1 i_2351 (.ZN (n_2183), .A (n_2215), .B (n_2184));
NAND2_X1 i_2350 (.ZN (n_2182), .A1 (B[23]), .A2 (A[11]));
XOR2_X1 i_2349 (.Z (n_2181), .A (n_2183), .B (n_2182));
XOR2_X1 i_2348 (.Z (n_2180), .A (n_2186), .B (n_2185));
XOR2_X1 i_2347 (.Z (n_2179), .A (n_2181), .B (n_2180));
AOI22_X1 i_2346 (.ZN (n_2178), .A1 (n_2181), .A2 (n_2180), .B1 (n_2194), .B2 (n_2179));
NAND2_X1 i_2345 (.ZN (n_2177), .A1 (B[13]), .A2 (A[21]));
NAND2_X1 i_2344 (.ZN (n_2176), .A1 (B[17]), .A2 (A[16]));
XNOR2_X1 i_2343 (.ZN (n_2175), .A (n_1965), .B (n_2176));
NAND2_X1 i_2342 (.ZN (n_2174), .A1 (B[15]), .A2 (A[18]));
OAI22_X1 i_2341 (.ZN (n_2173), .A1 (n_1965), .A2 (n_2176), .B1 (n_2175), .B2 (n_2174));
AOI22_X1 i_2340 (.ZN (n_2172), .A1 (B[13]), .A2 (A[20]), .B1 (B[12]), .B2 (A[21]));
INV_X1 i_2339 (.ZN (n_2154), .A (n_2172));
OAI21_X1 i_2338 (.ZN (n_2153), .A (n_2154), .B1 (n_1985), .B2 (n_2177));
OR2_X1 i_2337 (.ZN (n_2152), .A1 (n_559), .A2 (n_853));
OAI22_X1 i_2336 (.ZN (n_2151), .A1 (n_1985), .A2 (n_2177), .B1 (n_2153), .B2 (n_2152));
NAND2_X1 i_2335 (.ZN (n_2150), .A1 (n_2173), .A2 (n_2151));
OAI21_X1 i_2334 (.ZN (n_2149), .A (n_2150), .B1 (n_2173), .B2 (n_2151));
OAI21_X1 i_2333 (.ZN (n_2148), .A (n_2150), .B1 (n_2003), .B2 (n_2149));
OAI22_X1 i_2332 (.ZN (n_2147), .A1 (n_2215), .A2 (n_2184), .B1 (n_2183), .B2 (n_2182));
XOR2_X1 i_2331 (.Z (n_2146), .A (n_2148), .B (n_2147));
NOR2_X1 i_2330 (.ZN (n_2145), .A1 (n_559), .A2 (n_1792));
AND3_X1 i_2329 (.ZN (n_2143), .A1 (B[12]), .A2 (A[21]), .A3 (n_2145));
AOI22_X1 i_2328 (.ZN (n_2142), .A1 (B[12]), .A2 (A[23]), .B1 (B[14]), .B2 (A[21]));
NOR2_X1 i_2327 (.ZN (n_2137), .A1 (n_2143), .A2 (n_2142));
NOR2_X1 i_2326 (.ZN (n_2136), .A1 (n_229), .A2 (n_1881));
XOR2_X1 i_2325 (.Z (n_2135), .A (n_2137), .B (n_2136));
XOR2_X1 i_2324 (.Z (n_2134), .A (n_2146), .B (n_2135));
XNOR2_X1 i_2323 (.ZN (n_2133), .A (n_2178), .B (n_2134));
NAND2_X1 i_2322 (.ZN (n_2132), .A1 (B[21]), .A2 (A[10]));
XNOR2_X1 i_2321 (.ZN (n_2131), .A (n_1924), .B (n_2234));
NAND2_X1 i_2320 (.ZN (n_2130), .A1 (B[14]), .A2 (A[17]));
AOI21_X1 i_2319 (.ZN (n_2129), .A (n_2054), .B1 (n_2056), .B2 (n_2057));
OAI22_X1 i_2318 (.ZN (n_2128), .A1 (n_1924), .A2 (n_2234), .B1 (n_2131), .B2 (n_2130));
INV_X1 i_2317 (.ZN (n_2127), .A (n_2128));
NOR2_X1 i_2316 (.ZN (n_2126), .A1 (n_2129), .A2 (n_2127));
AOI21_X1 i_2315 (.ZN (n_2125), .A (n_2126), .B1 (n_2129), .B2 (n_2127));
OR2_X1 i_2314 (.ZN (n_2124), .A1 (n_1963), .A2 (n_1848));
AOI22_X1 i_2313 (.ZN (n_2123), .A1 (B[16]), .A2 (A[15]), .B1 (B[17]), .B2 (A[14]));
INV_X1 i_2312 (.ZN (n_2122), .A (n_2123));
NAND2_X1 i_2311 (.ZN (n_2119), .A1 (n_2124), .A2 (n_2122));
OAI21_X1 i_2310 (.ZN (n_2118), .A (n_2124), .B1 (n_1964), .B2 (n_2119));
OAI33_X1 i_2309 (.ZN (n_2117), .A1 (n_1235), .A2 (n_1368), .A3 (n_2132), .B1 (n_1979)
    , .B2 (n_339), .B3 (n_1533));
INV_X1 i_2308 (.ZN (n_2116), .A (n_2117));
AOI21_X1 i_2307 (.ZN (n_2115), .A (n_2126), .B1 (n_2125), .B2 (n_2118));
NOR2_X1 i_2306 (.ZN (n_2114), .A1 (n_2116), .A2 (n_2115));
AOI21_X1 i_2305 (.ZN (n_2111), .A (n_2114), .B1 (n_2116), .B2 (n_2115));
AOI21_X1 i_2304 (.ZN (n_2110), .A (n_2025), .B1 (n_2236), .B2 (n_2037));
NOR2_X1 i_2303 (.ZN (n_2109), .A1 (n_2243), .A2 (n_1792));
XOR2_X1 i_2302 (.Z (n_2108), .A (n_2110), .B (n_2109));
INV_X1 i_2301 (.ZN (n_2107), .A (n_2108));
NAND2_X1 i_2300 (.ZN (n_2088), .A1 (B[11]), .A2 (A[22]));
INV_X1 i_2299 (.ZN (n_2087), .A (n_2088));
OAI22_X1 i_2298 (.ZN (n_2086), .A1 (n_2107), .A2 (n_2088), .B1 (n_2108), .B2 (n_2087));
AOI21_X1 i_2297 (.ZN (n_2085), .A (n_2114), .B1 (n_2111), .B2 (n_2086));
XOR2_X1 i_2296 (.Z (n_2084), .A (n_1958), .B (n_2200));
XOR2_X1 i_2295 (.Z (n_2083), .A (n_2153), .B (n_2152));
NOR2_X1 i_2294 (.ZN (n_2082), .A1 (n_2084), .A2 (n_2083));
AOI21_X1 i_2293 (.ZN (n_2081), .A (n_2082), .B1 (n_2084), .B2 (n_2083));
XNOR2_X1 i_2292 (.ZN (n_2080), .A (n_2175), .B (n_2174));
XOR2_X1 i_2291 (.Z (n_2079), .A (n_2003), .B (n_2149));
AOI21_X1 i_2290 (.ZN (n_2078), .A (n_2082), .B1 (n_2081), .B2 (n_2080));
NOR2_X1 i_2289 (.ZN (n_2077), .A1 (n_2079), .A2 (n_2078));
AOI21_X1 i_2288 (.ZN (n_2076), .A (n_2077), .B1 (n_2079), .B2 (n_2078));
AOI21_X1 i_2287 (.ZN (n_2075), .A (n_2077), .B1 (n_2085), .B2 (n_2076));
XNOR2_X1 i_2286 (.ZN (n_2074), .A (n_2133), .B (n_2075));
AOI22_X1 i_2285 (.ZN (n_2073), .A1 (n_2071), .A2 (n_2072), .B1 (n_2069), .B2 (n_2070));
INV_X1 i_2284 (.ZN (n_2072), .A (n_2068));
XOR2_X1 i_2283 (.Z (n_2071), .A (n_2069), .B (n_2070));
XOR2_X1 i_2282 (.Z (n_2070), .A (n_1991), .B (n_2038));
XNOR2_X1 i_2281 (.ZN (n_2069), .A (n_1976), .B (n_1981));
OAI21_X1 i_2280 (.ZN (n_2068), .A (n_2063), .B1 (n_2064), .B2 (n_2067));
INV_X1 i_2279 (.ZN (n_2067), .A (n_2066));
AOI22_X1 i_2278 (.ZN (n_2066), .A1 (n_2065), .A2 (n_1796), .B1 (n_1811), .B2 (n_1797));
INV_X1 i_2277 (.ZN (n_2065), .A (n_1795));
OAI21_X1 i_2276 (.ZN (n_2064), .A (n_2063), .B1 (n_2062), .B2 (n_2061));
NAND2_X1 i_2275 (.ZN (n_2063), .A1 (n_2061), .A2 (n_2062));
AOI22_X1 i_2274 (.ZN (n_2062), .A1 (n_1842), .A2 (n_1833), .B1 (n_1832), .B2 (n_1813));
OAI21_X1 i_2273 (.ZN (n_2061), .A (n_2060), .B1 (n_2059), .B2 (n_2058));
NAND2_X1 i_2272 (.ZN (n_2060), .A1 (n_2058), .A2 (n_2059));
XNOR2_X1 i_2271 (.ZN (n_2059), .A (n_2053), .B (n_2041));
XOR2_X1 i_2270 (.Z (n_2058), .A (n_2056), .B (n_2057));
AND2_X1 i_2269 (.ZN (n_2057), .A1 (B[11]), .A2 (A[20]));
NOR2_X1 i_2268 (.ZN (n_2056), .A1 (n_2054), .A2 (n_2055));
AOI22_X1 i_2267 (.ZN (n_2055), .A1 (B[10]), .A2 (A[21]), .B1 (B[9]), .B2 (A[22]));
NOR2_X1 i_2266 (.ZN (n_2054), .A1 (n_1992), .A2 (n_1954));
AOI22_X1 i_2265 (.ZN (n_2053), .A1 (n_1850), .A2 (n_1853), .B1 (n_1849), .B2 (n_1843));
INV_X1 i_2264 (.ZN (n_2052), .A (n_2041));
OAI22_X1 i_2263 (.ZN (n_2041), .A1 (n_2039), .A2 (n_1934), .B1 (n_2040), .B2 (n_1726));
INV_X1 i_2262 (.ZN (n_2040), .A (n_1932));
INV_X1 i_2261 (.ZN (n_2039), .A (n_1933));
XNOR2_X1 i_2260 (.ZN (n_2038), .A (n_2037), .B (n_1992));
NOR2_X1 i_2259 (.ZN (n_2037), .A1 (n_2025), .A2 (n_2026));
AOI22_X1 i_2258 (.ZN (n_2026), .A1 (A[23]), .A2 (B[9]), .B1 (A[21]), .B2 (B[11]));
NOR2_X1 i_2257 (.ZN (n_2025), .A1 (n_2003), .A2 (n_1954));
NAND2_X1 i_2256 (.ZN (n_2003), .A1 (A[23]), .A2 (B[11]));
NAND2_X1 i_2255 (.ZN (n_1992), .A1 (B[10]), .A2 (A[22]));
XNOR2_X1 i_2254 (.ZN (n_1991), .A (n_1990), .B (n_1984));
XOR2_X1 i_2253 (.Z (n_1990), .A (n_1987), .B (n_1988));
NAND2_X1 i_2252 (.ZN (n_1988), .A1 (B[14]), .A2 (A[18]));
XNOR2_X1 i_2251 (.ZN (n_1987), .A (n_1985), .B (n_1986));
NAND2_X1 i_2250 (.ZN (n_1986), .A1 (B[13]), .A2 (A[19]));
NAND2_X1 i_2249 (.ZN (n_1985), .A1 (B[12]), .A2 (A[20]));
AOI22_X1 i_2248 (.ZN (n_1984), .A1 (n_1982), .A2 (n_1908), .B1 (n_1907), .B2 (n_1906));
INV_X1 i_2247 (.ZN (n_1982), .A (n_1909));
XNOR2_X1 i_2246 (.ZN (n_1981), .A (n_1979), .B (n_1980));
NAND2_X1 i_2245 (.ZN (n_1980), .A1 (B[23]), .A2 (A[9]));
XNOR2_X1 i_2244 (.ZN (n_1979), .A (n_1977), .B (n_1978));
NAND2_X1 i_2243 (.ZN (n_1978), .A1 (B[22]), .A2 (A[10]));
NAND2_X1 i_2242 (.ZN (n_1977), .A1 (B[21]), .A2 (A[11]));
XOR2_X1 i_2241 (.Z (n_1976), .A (n_1962), .B (n_1975));
XOR2_X1 i_2240 (.Z (n_1975), .A (n_1974), .B (n_1963));
NOR2_X1 i_2239 (.ZN (n_1974), .A1 (n_1966), .A2 (n_1967));
AOI22_X1 i_2238 (.ZN (n_1967), .A1 (B[15]), .A2 (A[17]), .B1 (B[16]), .B2 (A[16]));
NOR2_X1 i_2237 (.ZN (n_1966), .A1 (n_1964), .A2 (n_1965));
NAND2_X1 i_2236 (.ZN (n_1965), .A1 (A[17]), .A2 (B[16]));
NAND2_X1 i_2235 (.ZN (n_1964), .A1 (B[15]), .A2 (A[16]));
NAND2_X1 i_2234 (.ZN (n_1963), .A1 (B[17]), .A2 (A[15]));
XOR2_X1 i_2233 (.Z (n_1962), .A (n_1961), .B (n_1957));
NOR2_X1 i_2232 (.ZN (n_1961), .A1 (n_1959), .A2 (n_1960));
AOI22_X1 i_2231 (.ZN (n_1960), .A1 (B[19]), .A2 (A[13]), .B1 (B[20]), .B2 (A[12]));
NOR2_X1 i_2230 (.ZN (n_1959), .A1 (n_1958), .A2 (n_1929));
NAND2_X1 i_2229 (.ZN (n_1958), .A1 (A[13]), .A2 (B[20]));
NAND2_X1 i_2228 (.ZN (n_1957), .A1 (B[18]), .A2 (A[14]));
INV_X1 i_2227 (.ZN (n_1956), .A (n_1879));
INV_X1 i_2226 (.ZN (n_1955), .A (B[7]));
NAND2_X1 i_2225 (.ZN (n_1954), .A1 (B[9]), .A2 (A[21]));
NAND2_X1 i_2224 (.ZN (n_1953), .A1 (n_1886), .A2 (n_1885));
OAI21_X1 i_2223 (.ZN (n_1952), .A (n_1953), .B1 (n_1884), .B2 (n_1956));
XNOR2_X1 i_2222 (.ZN (n_1951), .A (n_1873), .B (n_1954));
NAND2_X1 i_2221 (.ZN (n_1941), .A1 (B[11]), .A2 (A[19]));
XOR2_X1 i_2220 (.Z (n_1936), .A (n_1951), .B (n_1941));
XOR2_X1 i_2219 (.Z (n_1935), .A (n_1952), .B (n_1936));
AOI21_X1 i_2218 (.ZN (n_1934), .A (n_1725), .B1 (n_1723), .B2 (n_1722));
NOR2_X1 i_2217 (.ZN (n_1933), .A1 (n_1955), .A2 (n_1792));
XNOR2_X1 i_2216 (.ZN (n_1932), .A (n_1934), .B (n_1933));
XNOR2_X1 i_2215 (.ZN (n_1931), .A (n_1726), .B (n_1932));
AOI22_X1 i_2214 (.ZN (n_1930), .A1 (n_1952), .A2 (n_1936), .B1 (n_1935), .B2 (n_1931));
NAND2_X1 i_2213 (.ZN (n_1929), .A1 (B[19]), .A2 (A[12]));
NOR3_X1 i_2212 (.ZN (n_1928), .A1 (n_1235), .A2 (n_1929), .A3 (n_1532));
AOI22_X1 i_2211 (.ZN (n_1927), .A1 (B[19]), .A2 (A[11]), .B1 (B[18]), .B2 (A[12]));
NOR2_X1 i_2210 (.ZN (n_1926), .A1 (n_1928), .A2 (n_1927));
NOR2_X1 i_2209 (.ZN (n_1925), .A1 (n_1339), .A2 (n_856));
NAND2_X1 i_2208 (.ZN (n_1924), .A1 (B[13]), .A2 (A[18]));
NOR2_X1 i_2207 (.ZN (n_1923), .A1 (n_1852), .A2 (n_1924));
AOI22_X1 i_2206 (.ZN (n_1922), .A1 (B[13]), .A2 (A[17]), .B1 (B[12]), .B2 (A[18]));
OR2_X1 i_2205 (.ZN (n_1921), .A1 (n_1923), .A2 (n_1922));
OR2_X1 i_2204 (.ZN (n_1920), .A1 (n_559), .A2 (n_1305));
NOR2_X1 i_2203 (.ZN (n_1918), .A1 (n_1921), .A2 (n_1920));
AOI21_X1 i_2202 (.ZN (n_1917), .A (n_1918), .B1 (n_1921), .B2 (n_1920));
XOR2_X1 i_2201 (.Z (n_1916), .A (n_1926), .B (n_1925));
NOR2_X1 i_2200 (.ZN (n_1915), .A1 (n_1917), .A2 (n_1916));
AOI21_X1 i_2199 (.ZN (n_1914), .A (n_1915), .B1 (n_1917), .B2 (n_1916));
NAND2_X1 i_2198 (.ZN (n_1913), .A1 (B[17]), .A2 (A[13]));
XNOR2_X1 i_2197 (.ZN (n_1912), .A (n_1848), .B (n_1913));
NAND2_X1 i_2196 (.ZN (n_1911), .A1 (B[15]), .A2 (A[15]));
XNOR2_X1 i_2195 (.ZN (n_1910), .A (n_1912), .B (n_1911));
NOR2_X1 i_2194 (.ZN (n_1909), .A1 (n_1923), .A2 (n_1918));
NOR2_X1 i_2193 (.ZN (n_1908), .A1 (n_1792), .A2 (n_425));
XNOR2_X1 i_2192 (.ZN (n_1907), .A (n_1909), .B (n_1908));
OAI22_X1 i_2191 (.ZN (n_1906), .A1 (n_1873), .A2 (n_1954), .B1 (n_1951), .B2 (n_1941));
AOI21_X1 i_2190 (.ZN (n_1905), .A (n_1915), .B1 (n_1914), .B2 (n_1910));
XOR2_X1 i_2189 (.Z (n_1897), .A (n_1907), .B (n_1906));
NOR2_X1 i_2188 (.ZN (n_1896), .A1 (n_1905), .A2 (n_1897));
AOI21_X1 i_2187 (.ZN (n_1895), .A (n_1896), .B1 (n_1905), .B2 (n_1897));
AOI21_X1 i_2186 (.ZN (n_1894), .A (n_1896), .B1 (n_1930), .B2 (n_1895));
INV_X1 i_2185 (.ZN (n_1893), .A (n_1883));
OAI21_X1 i_2184 (.ZN (n_1892), .A (n_1891), .B1 (n_1888), .B2 (n_1887));
NAND2_X1 i_2183 (.ZN (n_1891), .A1 (n_1889), .A2 (n_1890));
AOI22_X1 i_2182 (.ZN (n_1890), .A1 (n_1709), .A2 (n_1716), .B1 (n_1703), .B2 (n_1708));
XOR2_X1 i_2181 (.Z (n_1889), .A (n_1887), .B (n_1888));
XNOR2_X1 i_2180 (.ZN (n_1888), .A (n_1828), .B (n_1824));
XNOR2_X1 i_2179 (.ZN (n_1887), .A (n_1886), .B (n_1885));
XNOR2_X1 i_2178 (.ZN (n_1886), .A (n_1879), .B (n_1884));
OAI21_X1 i_2177 (.ZN (n_1885), .A (n_1699), .B1 (n_1701), .B2 (n_1702));
OAI21_X1 i_2176 (.ZN (n_1884), .A (n_1880), .B1 (n_1883), .B2 (n_1882));
NOR3_X1 i_2175 (.ZN (n_1883), .A1 (n_1783), .A2 (n_425), .A3 (n_1322));
NOR2_X1 i_2174 (.ZN (n_1882), .A1 (n_1881), .A2 (n_169));
INV_X1 i_2173 (.ZN (n_1881), .A (A[22]));
OAI21_X1 i_2172 (.ZN (n_1880), .A (n_1783), .B1 (n_425), .B2 (n_1322));
OAI22_X1 i_2171 (.ZN (n_1879), .A1 (n_1877), .A2 (n_1878), .B1 (n_1876), .B2 (n_1874));
NAND2_X1 i_2170 (.ZN (n_1878), .A1 (B[11]), .A2 (A[17]));
XNOR2_X1 i_2169 (.ZN (n_1877), .A (n_1876), .B (n_1874));
NAND2_X1 i_2168 (.ZN (n_1876), .A1 (B[10]), .A2 (A[18]));
INV_X1 i_2167 (.ZN (n_1875), .A (n_1568));
NAND2_X1 i_2166 (.ZN (n_1874), .A1 (B[9]), .A2 (A[19]));
NAND2_X1 i_2165 (.ZN (n_1873), .A1 (B[10]), .A2 (A[20]));
AND2_X1 i_2164 (.ZN (n_1872), .A1 (B[9]), .A2 (A[20]));
AND2_X1 i_2163 (.ZN (n_1871), .A1 (B[10]), .A2 (A[19]));
NAND2_X1 i_2162 (.ZN (n_1870), .A1 (n_1872), .A2 (n_1871));
OAI21_X1 i_2161 (.ZN (n_1869), .A (n_1870), .B1 (n_1872), .B2 (n_1871));
NAND2_X1 i_2160 (.ZN (n_1868), .A1 (B[11]), .A2 (A[18]));
OAI21_X1 i_2159 (.ZN (n_1853), .A (n_1870), .B1 (n_1869), .B2 (n_1868));
NAND2_X1 i_2158 (.ZN (n_1852), .A1 (B[12]), .A2 (A[17]));
XNOR2_X1 i_2157 (.ZN (n_1851), .A (n_1698), .B (n_1852));
OAI33_X1 i_2156 (.ZN (n_1850), .A1 (n_559), .A2 (n_558), .A3 (n_1851), .B1 (n_229)
    , .B2 (n_1305), .B3 (n_1852));
XOR2_X1 i_2155 (.Z (n_1849), .A (n_1853), .B (n_1850));
NAND2_X1 i_2154 (.ZN (n_1848), .A1 (B[16]), .A2 (A[14]));
AOI22_X1 i_2153 (.ZN (n_1847), .A1 (B[16]), .A2 (A[13]), .B1 (B[15]), .B2 (A[14]));
INV_X1 i_2152 (.ZN (n_1846), .A (n_1847));
OAI21_X1 i_2151 (.ZN (n_1845), .A (n_1846), .B1 (n_1707), .B2 (n_1848));
NAND2_X1 i_2150 (.ZN (n_1844), .A1 (B[17]), .A2 (A[12]));
OAI22_X1 i_2149 (.ZN (n_1843), .A1 (n_1707), .A2 (n_1848), .B1 (n_1845), .B2 (n_1844));
XOR2_X1 i_2148 (.Z (n_1842), .A (n_1849), .B (n_1843));
NAND2_X1 i_2147 (.ZN (n_1841), .A1 (B[23]), .A2 (A[7]));
NAND2_X1 i_2146 (.ZN (n_1840), .A1 (B[22]), .A2 (A[9]));
NOR3_X1 i_2145 (.ZN (n_1839), .A1 (n_458), .A2 (n_1840), .A3 (n_1367));
INV_X1 i_2144 (.ZN (n_1838), .A (n_1839));
AOI22_X1 i_2143 (.ZN (n_1837), .A1 (B[21]), .A2 (A[9]), .B1 (B[22]), .B2 (A[8]));
NOR2_X1 i_2142 (.ZN (n_1834), .A1 (n_1839), .A2 (n_1837));
XNOR2_X1 i_2141 (.ZN (n_1833), .A (n_1841), .B (n_1834));
XOR2_X1 i_2140 (.Z (n_1832), .A (n_1842), .B (n_1833));
OAI22_X1 i_2139 (.ZN (n_1831), .A1 (n_1707), .A2 (n_1706), .B1 (n_1704), .B2 (n_1705));
INV_X1 i_2138 (.ZN (n_1830), .A (n_1831));
AOI21_X1 i_2137 (.ZN (n_1829), .A (n_1712), .B1 (n_1714), .B2 (n_1715));
XNOR2_X1 i_2136 (.ZN (n_1828), .A (n_1830), .B (n_1829));
NOR2_X1 i_2135 (.ZN (n_1827), .A1 (n_1460), .A2 (n_1567));
AOI22_X1 i_2134 (.ZN (n_1826), .A1 (B[23]), .A2 (A[5]), .B1 (B[22]), .B2 (A[6]));
NOR2_X1 i_2133 (.ZN (n_1825), .A1 (n_1827), .A2 (n_1826));
AOI21_X1 i_2132 (.ZN (n_1824), .A (n_1827), .B1 (n_1573), .B2 (n_1825));
OAI22_X1 i_2131 (.ZN (n_1823), .A1 (n_1830), .A2 (n_1829), .B1 (n_1828), .B2 (n_1824));
AOI21_X1 i_2130 (.ZN (n_1822), .A (n_1875), .B1 (n_1567), .B2 (n_1569));
INV_X1 i_2129 (.ZN (n_1821), .A (n_1822));
AOI21_X1 i_2128 (.ZN (n_1815), .A (n_1559), .B1 (n_1558), .B2 (n_1557));
XOR2_X1 i_2127 (.Z (n_1814), .A (n_1822), .B (n_1815));
XOR2_X1 i_2126 (.Z (n_1813), .A (n_1823), .B (n_1814));
XOR2_X1 i_2125 (.Z (n_1812), .A (n_1832), .B (n_1813));
AOI22_X1 i_2124 (.ZN (n_1811), .A1 (n_1720), .A2 (n_1757), .B1 (n_1728), .B2 (n_1721));
XOR2_X1 i_2123 (.Z (n_1810), .A (n_1869), .B (n_1868));
NAND2_X1 i_2122 (.ZN (n_1809), .A1 (B[14]), .A2 (A[15]));
XOR2_X1 i_2121 (.Z (n_1808), .A (n_1851), .B (n_1809));
NOR2_X1 i_2120 (.ZN (n_1807), .A1 (n_1810), .A2 (n_1808));
AOI21_X1 i_2119 (.ZN (n_1806), .A (n_1807), .B1 (n_1810), .B2 (n_1808));
XNOR2_X1 i_2118 (.ZN (n_1805), .A (n_1845), .B (n_1844));
AOI21_X1 i_2117 (.ZN (n_1797), .A (n_1807), .B1 (n_1806), .B2 (n_1805));
XOR2_X1 i_2116 (.Z (n_1796), .A (n_1811), .B (n_1797));
AOI22_X1 i_2115 (.ZN (n_1795), .A1 (n_1574), .A2 (n_1553), .B1 (n_1563), .B2 (n_1554));
XNOR2_X1 i_2114 (.ZN (n_1794), .A (n_1796), .B (n_1795));
XOR2_X1 i_2113 (.Z (n_1793), .A (n_1812), .B (n_1794));
INV_X1 i_2112 (.ZN (n_1792), .A (A[23]));
INV_X1 i_2111 (.ZN (n_1791), .A (n_1607));
INV_X1 i_2110 (.ZN (n_1790), .A (n_1590));
NAND2_X1 i_2109 (.ZN (n_1789), .A1 (B[11]), .A2 (A[16]));
XNOR2_X1 i_2108 (.ZN (n_1788), .A (n_1630), .B (n_1789));
NAND2_X1 i_2107 (.ZN (n_1787), .A1 (B[9]), .A2 (A[18]));
NOR2_X1 i_2106 (.ZN (n_1786), .A1 (n_1792), .A2 (n_1029));
OAI22_X1 i_2105 (.ZN (n_1785), .A1 (n_1630), .A2 (n_1789), .B1 (n_1788), .B2 (n_1787));
XOR2_X1 i_2104 (.Z (n_1784), .A (n_1786), .B (n_1785));
NAND2_X1 i_2103 (.ZN (n_1783), .A1 (B[7]), .A2 (A[21]));
NOR2_X1 i_2102 (.ZN (n_1782), .A1 (n_1635), .A2 (n_1783));
AOI22_X1 i_2101 (.ZN (n_1763), .A1 (B[6]), .A2 (A[21]), .B1 (B[7]), .B2 (A[20]));
NOR2_X1 i_2100 (.ZN (n_1762), .A1 (n_1782), .A2 (n_1763));
OAI22_X1 i_2099 (.ZN (n_1761), .A1 (n_1635), .A2 (n_1783), .B1 (n_1648), .B2 (n_1763));
INV_X1 i_2098 (.ZN (n_1760), .A (n_1761));
AOI22_X1 i_2097 (.ZN (n_1757), .A1 (n_1786), .A2 (n_1785), .B1 (n_1784), .B2 (n_1761));
NOR2_X1 i_2096 (.ZN (n_1755), .A1 (n_1603), .A2 (n_1704));
AOI22_X1 i_2095 (.ZN (n_1754), .A1 (B[15]), .A2 (A[12]), .B1 (B[16]), .B2 (A[11]));
NOR2_X1 i_2094 (.ZN (n_1746), .A1 (n_1755), .A2 (n_1754));
NAND2_X1 i_2093 (.ZN (n_1745), .A1 (n_1791), .A2 (n_1746));
NOR2_X1 i_2092 (.ZN (n_1744), .A1 (n_1676), .A2 (n_558));
NOR2_X1 i_2091 (.ZN (n_1743), .A1 (n_229), .A2 (n_557));
NAND2_X1 i_2090 (.ZN (n_1740), .A1 (n_1744), .A2 (n_1743));
OAI21_X1 i_2089 (.ZN (n_1739), .A (n_1740), .B1 (n_1744), .B2 (n_1743));
NAND2_X1 i_2088 (.ZN (n_1738), .A1 (B[14]), .A2 (A[13]));
OAI21_X1 i_2087 (.ZN (n_1737), .A (n_1745), .B1 (n_1603), .B2 (n_1704));
OAI21_X1 i_2086 (.ZN (n_1736), .A (n_1740), .B1 (n_1739), .B2 (n_1738));
XOR2_X1 i_2085 (.Z (n_1734), .A (n_1737), .B (n_1736));
NOR2_X1 i_2084 (.ZN (n_1733), .A1 (n_556), .A2 (n_856));
NAND2_X1 i_2083 (.ZN (n_1732), .A1 (n_1790), .A2 (n_1733));
OAI21_X1 i_2082 (.ZN (n_1731), .A (n_1732), .B1 (n_1790), .B2 (n_1733));
OAI21_X1 i_2081 (.ZN (n_1730), .A (n_1732), .B1 (n_1710), .B2 (n_1731));
AOI22_X1 i_2080 (.ZN (n_1728), .A1 (n_1737), .A2 (n_1736), .B1 (n_1734), .B2 (n_1730));
NAND2_X1 i_2079 (.ZN (n_1726), .A1 (B[8]), .A2 (A[22]));
NOR2_X1 i_2078 (.ZN (n_1725), .A1 (n_1783), .A2 (n_1726));
AOI22_X1 i_2077 (.ZN (n_1724), .A1 (B[7]), .A2 (A[22]), .B1 (B[8]), .B2 (A[21]));
NOR2_X1 i_2076 (.ZN (n_1723), .A1 (n_1725), .A2 (n_1724));
NOR2_X1 i_2075 (.ZN (n_1722), .A1 (n_1792), .A2 (n_169));
XNOR2_X1 i_2074 (.ZN (n_1721), .A (n_1723), .B (n_1722));
XOR2_X1 i_2073 (.Z (n_1720), .A (n_1728), .B (n_1721));
XOR2_X1 i_2072 (.Z (n_1719), .A (n_1757), .B (n_1720));
AOI21_X1 i_2071 (.ZN (n_1718), .A (n_1661), .B1 (n_1717), .B2 (n_1662));
XNOR2_X1 i_2070 (.ZN (n_1717), .A (n_1709), .B (n_1716));
XNOR2_X1 i_2069 (.ZN (n_1716), .A (n_1714), .B (n_1715));
NOR2_X1 i_2068 (.ZN (n_1715), .A1 (n_458), .A2 (n_856));
NOR2_X1 i_2067 (.ZN (n_1714), .A1 (n_1712), .A2 (n_1713));
AOI22_X1 i_2066 (.ZN (n_1713), .A1 (B[19]), .A2 (A[9]), .B1 (B[18]), .B2 (A[10]));
NOR3_X1 i_2065 (.ZN (n_1712), .A1 (n_1710), .A2 (n_1711), .A3 (n_1339));
INV_X1 i_2064 (.ZN (n_1711), .A (B[19]));
NAND2_X1 i_2063 (.ZN (n_1710), .A1 (A[9]), .A2 (B[18]));
XOR2_X1 i_2062 (.Z (n_1709), .A (n_1708), .B (n_1703));
XNOR2_X1 i_2061 (.ZN (n_1708), .A (n_1706), .B (n_1707));
NAND2_X1 i_2060 (.ZN (n_1707), .A1 (B[15]), .A2 (A[13]));
XNOR2_X1 i_2059 (.ZN (n_1706), .A (n_1704), .B (n_1705));
NAND2_X1 i_2058 (.ZN (n_1705), .A1 (B[17]), .A2 (A[11]));
NAND2_X1 i_2057 (.ZN (n_1704), .A1 (B[16]), .A2 (A[12]));
XNOR2_X1 i_2056 (.ZN (n_1703), .A (n_1701), .B (n_1702));
NAND2_X1 i_2055 (.ZN (n_1702), .A1 (B[14]), .A2 (A[14]));
NAND2_X1 i_2054 (.ZN (n_1701), .A1 (n_1699), .A2 (n_1700));
OAI22_X1 i_2053 (.ZN (n_1700), .A1 (n_1676), .A2 (n_1305), .B1 (n_558), .B2 (n_229));
OR3_X1 i_2052 (.ZN (n_1699), .A1 (n_1698), .A2 (n_1676), .A3 (n_558));
NAND2_X1 i_2051 (.ZN (n_1698), .A1 (B[13]), .A2 (A[16]));
INV_X1 i_2050 (.ZN (n_1676), .A (B[12]));
AOI21_X1 i_2049 (.ZN (n_1662), .A (n_1661), .B1 (n_1659), .B2 (n_1660));
NOR2_X1 i_2048 (.ZN (n_1661), .A1 (n_1659), .A2 (n_1660));
XOR2_X1 i_2047 (.Z (n_1660), .A (n_1608), .B (n_1575));
AOI22_X1 i_2046 (.ZN (n_1659), .A1 (n_1655), .A2 (n_1658), .B1 (n_1650), .B2 (n_1654));
XNOR2_X1 i_2045 (.ZN (n_1658), .A (n_1620), .B (n_1614));
XOR2_X1 i_2044 (.Z (n_1655), .A (n_1650), .B (n_1654));
OAI22_X1 i_2043 (.ZN (n_1654), .A1 (n_1652), .A2 (n_1366), .B1 (n_1653), .B2 (n_1447));
INV_X1 i_2042 (.ZN (n_1653), .A (n_1374));
INV_X1 i_2041 (.ZN (n_1652), .A (n_1373));
XNOR2_X1 i_2040 (.ZN (n_1650), .A (n_1579), .B (n_1577));
INV_X1 i_2039 (.ZN (n_1649), .A (n_1460));
NAND2_X1 i_2038 (.ZN (n_1648), .A1 (B[8]), .A2 (A[19]));
NOR2_X1 i_2037 (.ZN (n_1647), .A1 (n_1375), .A2 (n_1648));
AOI22_X1 i_2036 (.ZN (n_1640), .A1 (B[8]), .A2 (A[18]), .B1 (B[7]), .B2 (A[19]));
NOR2_X1 i_2035 (.ZN (n_1636), .A1 (n_1647), .A2 (n_1640));
NAND2_X1 i_2034 (.ZN (n_1635), .A1 (B[6]), .A2 (A[20]));
INV_X1 i_2033 (.ZN (n_1634), .A (n_1635));
NAND2_X1 i_2032 (.ZN (n_1631), .A1 (B[9]), .A2 (A[16]));
NAND2_X1 i_2031 (.ZN (n_1630), .A1 (B[10]), .A2 (A[17]));
NOR2_X1 i_2030 (.ZN (n_1629), .A1 (n_1631), .A2 (n_1630));
AOI22_X1 i_2029 (.ZN (n_1628), .A1 (B[10]), .A2 (A[16]), .B1 (B[9]), .B2 (A[17]));
NOR2_X1 i_2028 (.ZN (n_1627), .A1 (n_1629), .A2 (n_1628));
AND2_X1 i_2027 (.ZN (n_1626), .A1 (B[11]), .A2 (A[15]));
AOI21_X1 i_2026 (.ZN (n_1624), .A (n_1647), .B1 (n_1636), .B2 (n_1634));
AOI21_X1 i_2025 (.ZN (n_1623), .A (n_1629), .B1 (n_1627), .B2 (n_1626));
NOR2_X1 i_2024 (.ZN (n_1622), .A1 (n_1624), .A2 (n_1623));
AOI21_X1 i_2023 (.ZN (n_1621), .A (n_1622), .B1 (n_1624), .B2 (n_1623));
INV_X1 i_2022 (.ZN (n_1620), .A (n_1621));
NAND2_X1 i_2021 (.ZN (n_1617), .A1 (B[12]), .A2 (A[14]));
XNOR2_X1 i_2020 (.ZN (n_1616), .A (n_1529), .B (n_1617));
NAND2_X1 i_2019 (.ZN (n_1615), .A1 (B[14]), .A2 (A[12]));
OAI22_X1 i_2018 (.ZN (n_1614), .A1 (n_1529), .A2 (n_1617), .B1 (n_1616), .B2 (n_1615));
NOR2_X1 i_2017 (.ZN (n_1613), .A1 (n_170), .A2 (n_1367));
XOR2_X1 i_2016 (.Z (n_1612), .A (n_1649), .B (n_1613));
NOR2_X1 i_2015 (.ZN (n_1611), .A1 (n_422), .A2 (n_1533));
AOI21_X1 i_2014 (.ZN (n_1610), .A (n_1622), .B1 (n_1621), .B2 (n_1614));
AOI22_X1 i_2013 (.ZN (n_1609), .A1 (n_1649), .A2 (n_1613), .B1 (n_1612), .B2 (n_1611));
XOR2_X1 i_2012 (.Z (n_1608), .A (n_1610), .B (n_1609));
NAND2_X1 i_2011 (.ZN (n_1607), .A1 (B[17]), .A2 (A[10]));
NOR2_X1 i_2010 (.ZN (n_1606), .A1 (n_1524), .A2 (n_1607));
AOI22_X1 i_2009 (.ZN (n_1605), .A1 (B[17]), .A2 (A[9]), .B1 (B[16]), .B2 (A[10]));
NOR2_X1 i_2008 (.ZN (n_1604), .A1 (n_1606), .A2 (n_1605));
NAND2_X1 i_2007 (.ZN (n_1603), .A1 (B[15]), .A2 (A[11]));
INV_X1 i_2006 (.ZN (n_1602), .A (n_1603));
NAND2_X1 i_2005 (.ZN (n_1601), .A1 (n_1604), .A2 (n_1602));
NAND2_X1 i_2004 (.ZN (n_1590), .A1 (B[19]), .A2 (A[8]));
NOR2_X1 i_2003 (.ZN (n_1589), .A1 (n_1504), .A2 (n_1590));
AOI22_X1 i_2002 (.ZN (n_1588), .A1 (B[19]), .A2 (A[7]), .B1 (B[18]), .B2 (A[8]));
NOR2_X1 i_2001 (.ZN (n_1587), .A1 (n_1589), .A2 (n_1588));
OAI21_X1 i_2000 (.ZN (n_1586), .A (n_1601), .B1 (n_1524), .B2 (n_1607));
OAI22_X1 i_1999 (.ZN (n_1580), .A1 (n_1504), .A2 (n_1590), .B1 (n_1508), .B2 (n_1588));
XOR2_X1 i_1998 (.Z (n_1579), .A (n_1586), .B (n_1580));
AOI21_X1 i_1997 (.ZN (n_1577), .A (n_1459), .B1 (n_1455), .B2 (n_1454));
INV_X1 i_1996 (.ZN (n_1576), .A (n_1577));
AOI22_X1 i_1995 (.ZN (n_1575), .A1 (n_1586), .A2 (n_1580), .B1 (n_1579), .B2 (n_1576));
AOI22_X1 i_1994 (.ZN (n_1574), .A1 (n_1610), .A2 (n_1609), .B1 (n_1608), .B2 (n_1575));
NOR2_X1 i_1993 (.ZN (n_1573), .A1 (n_1367), .A2 (n_556));
NAND3_X1 i_1992 (.ZN (n_1569), .A1 (A[8]), .A2 (n_1573), .A3 (B[22]));
OAI22_X1 i_1991 (.ZN (n_1568), .A1 (n_1367), .A2 (n_458), .B1 (n_556), .B2 (n_1368));
NAND2_X1 i_1990 (.ZN (n_1567), .A1 (B[23]), .A2 (A[6]));
NAND2_X1 i_1989 (.ZN (n_1566), .A1 (n_1569), .A2 (n_1568));
XOR2_X1 i_1988 (.Z (n_1563), .A (n_1567), .B (n_1566));
NAND2_X1 i_1987 (.ZN (n_1562), .A1 (B[18]), .A2 (A[11]));
NAND2_X1 i_1986 (.ZN (n_1561), .A1 (B[19]), .A2 (A[10]));
NAND2_X1 i_1985 (.ZN (n_1560), .A1 (n_1562), .A2 (n_1561));
INV_X1 i_1984 (.ZN (n_1559), .A (n_1560));
OR2_X1 i_1983 (.ZN (n_1558), .A1 (n_1562), .A2 (n_1561));
NAND2_X1 i_1982 (.ZN (n_1557), .A1 (B[20]), .A2 (A[9]));
NAND2_X1 i_1981 (.ZN (n_1555), .A1 (n_1560), .A2 (n_1558));
XOR2_X1 i_1980 (.Z (n_1554), .A (n_1557), .B (n_1555));
XOR2_X1 i_1979 (.Z (n_1553), .A (n_1563), .B (n_1554));
XNOR2_X1 i_1978 (.ZN (n_1535), .A (n_1574), .B (n_1553));
INV_X1 i_1977 (.ZN (n_1534), .A (A[1]));
INV_X1 i_1976 (.ZN (n_1533), .A (B[23]));
INV_X1 i_1975 (.ZN (n_1532), .A (B[18]));
INV_X1 i_1974 (.ZN (n_1531), .A (n_1222));
INV_X1 i_1973 (.ZN (n_1530), .A (n_1262));
NAND2_X1 i_1972 (.ZN (n_1529), .A1 (A[13]), .A2 (B[13]));
AOI22_X1 i_1971 (.ZN (n_1528), .A1 (A[13]), .A2 (B[12]), .B1 (A[12]), .B2 (B[13]));
INV_X1 i_1970 (.ZN (n_1527), .A (n_1528));
OAI21_X1 i_1969 (.ZN (n_1526), .A (n_1527), .B1 (n_1343), .B2 (n_1529));
OAI22_X1 i_1968 (.ZN (n_1525), .A1 (n_1343), .A2 (n_1529), .B1 (n_1341), .B2 (n_1526));
NAND2_X1 i_1967 (.ZN (n_1524), .A1 (A[9]), .A2 (B[16]));
NAND2_X1 i_1966 (.ZN (n_1523), .A1 (A[10]), .A2 (B[15]));
XNOR2_X1 i_1965 (.ZN (n_1522), .A (n_1524), .B (n_1523));
OAI33_X1 i_1964 (.ZN (n_1521), .A1 (n_458), .A2 (n_1232), .A3 (n_1522), .B1 (n_1363)
    , .B2 (n_1339), .B3 (n_592));
XOR2_X1 i_1963 (.Z (n_1509), .A (n_1525), .B (n_1521));
NAND2_X1 i_1962 (.ZN (n_1508), .A1 (A[6]), .A2 (B[20]));
AOI22_X1 i_1961 (.ZN (n_1507), .A1 (A[5]), .A2 (B[20]), .B1 (A[6]), .B2 (B[19]));
INV_X1 i_1960 (.ZN (n_1506), .A (n_1507));
OAI21_X1 i_1959 (.ZN (n_1505), .A (n_1506), .B1 (n_1205), .B2 (n_1508));
NAND2_X1 i_1958 (.ZN (n_1504), .A1 (A[7]), .A2 (B[18]));
OAI22_X1 i_1957 (.ZN (n_1503), .A1 (n_1205), .A2 (n_1508), .B1 (n_1505), .B2 (n_1504));
XOR2_X1 i_1956 (.Z (n_1502), .A (n_1509), .B (n_1503));
AOI22_X1 i_1955 (.ZN (n_1501), .A1 (n_1212), .A2 (n_1198), .B1 (n_1531), .B2 (n_1213));
OAI22_X1 i_1954 (.ZN (n_1485), .A1 (n_99), .A2 (n_1367), .B1 (n_33), .B2 (n_1368));
NAND3_X1 i_1953 (.ZN (n_1484), .A1 (A[3]), .A2 (n_1530), .A3 (B[22]));
INV_X1 i_1952 (.ZN (n_1483), .A (n_1484));
NOR2_X1 i_1951 (.ZN (n_1482), .A1 (n_1534), .A2 (n_1533));
OAI21_X1 i_1950 (.ZN (n_1481), .A (n_1205), .B1 (n_1532), .B2 (n_170));
NOR3_X1 i_1949 (.ZN (n_1480), .A1 (n_1205), .A2 (n_170), .A3 (n_1532));
INV_X1 i_1948 (.ZN (n_1479), .A (n_1480));
NOR2_X1 i_1947 (.ZN (n_1478), .A1 (n_422), .A2 (n_856));
OAI21_X1 i_1946 (.ZN (n_1477), .A (n_1485), .B1 (n_1483), .B2 (n_1482));
OAI21_X1 i_1945 (.ZN (n_1476), .A (n_1481), .B1 (n_1480), .B2 (n_1478));
XNOR2_X1 i_1944 (.ZN (n_1461), .A (n_1477), .B (n_1476));
NAND2_X1 i_1943 (.ZN (n_1460), .A1 (A[5]), .A2 (B[22]));
NOR3_X1 i_1942 (.ZN (n_1459), .A1 (n_422), .A2 (n_1460), .A3 (n_1367));
AOI22_X1 i_1941 (.ZN (n_1456), .A1 (A[5]), .A2 (B[21]), .B1 (A[4]), .B2 (B[22]));
NOR2_X1 i_1940 (.ZN (n_1455), .A1 (n_1459), .A2 (n_1456));
NOR2_X1 i_1939 (.ZN (n_1454), .A1 (n_1533), .A2 (n_99));
OAI22_X1 i_1938 (.ZN (n_1453), .A1 (n_1477), .A2 (n_1476), .B1 (n_1501), .B2 (n_1461));
XOR2_X1 i_1937 (.Z (n_1452), .A (n_1455), .B (n_1454));
XOR2_X1 i_1936 (.Z (n_1450), .A (n_1453), .B (n_1452));
AOI22_X1 i_1935 (.ZN (n_1449), .A1 (n_1453), .A2 (n_1452), .B1 (n_1502), .B2 (n_1450));
INV_X1 i_1934 (.ZN (n_1448), .A (n_1449));
INV_X1 i_1933 (.ZN (n_1447), .A (n_1410));
AOI22_X1 i_1932 (.ZN (n_1444), .A1 (n_1413), .A2 (n_1443), .B1 (n_1411), .B2 (n_1412));
AOI22_X1 i_1931 (.ZN (n_1443), .A1 (n_1423), .A2 (n_1442), .B1 (n_1421), .B2 (n_1422));
OAI21_X1 i_1930 (.ZN (n_1442), .A (n_1441), .B1 (n_1425), .B2 (n_1424));
NAND2_X1 i_1929 (.ZN (n_1441), .A1 (n_1426), .A2 (n_1436));
XNOR2_X1 i_1928 (.ZN (n_1436), .A (n_1332), .B (n_1334));
XOR2_X1 i_1927 (.Z (n_1426), .A (n_1424), .B (n_1425));
XOR2_X1 i_1926 (.Z (n_1425), .A (n_1404), .B (n_1405));
XOR2_X1 i_1925 (.Z (n_1424), .A (n_1382), .B (n_1383));
XOR2_X1 i_1924 (.Z (n_1423), .A (n_1421), .B (n_1422));
XNOR2_X1 i_1923 (.ZN (n_1422), .A (n_1409), .B (n_1328));
AOI22_X1 i_1922 (.ZN (n_1421), .A1 (n_1418), .A2 (n_1420), .B1 (n_1414), .B2 (n_1415));
XOR2_X1 i_1921 (.Z (n_1420), .A (n_1364), .B (n_1419));
NAND2_X1 i_1920 (.ZN (n_1419), .A1 (A[7]), .A2 (B[17]));
XOR2_X1 i_1919 (.Z (n_1418), .A (n_1414), .B (n_1415));
XOR2_X1 i_1918 (.Z (n_1415), .A (n_1348), .B (n_1343));
XOR2_X1 i_1917 (.Z (n_1414), .A (n_1360), .B (n_1164));
XOR2_X1 i_1916 (.Z (n_1413), .A (n_1411), .B (n_1412));
OAI22_X1 i_1915 (.ZN (n_1412), .A1 (n_1326), .A2 (n_1338), .B1 (n_1324), .B2 (n_1325));
XOR2_X1 i_1914 (.Z (n_1411), .A (n_1374), .B (n_1410));
OAI22_X1 i_1913 (.ZN (n_1410), .A1 (n_1409), .A2 (n_1328), .B1 (n_1384), .B2 (n_1406));
XNOR2_X1 i_1912 (.ZN (n_1409), .A (n_1384), .B (n_1406));
AOI21_X1 i_1911 (.ZN (n_1406), .A (n_1402), .B1 (n_1404), .B2 (n_1405));
AND2_X1 i_1910 (.ZN (n_1405), .A1 (A[16]), .A2 (B[8]));
NOR2_X1 i_1909 (.ZN (n_1404), .A1 (n_1402), .A2 (n_1403));
AOI22_X1 i_1908 (.ZN (n_1403), .A1 (A[17]), .A2 (B[7]), .B1 (A[18]), .B2 (B[6]));
NOR2_X1 i_1907 (.ZN (n_1402), .A1 (n_1375), .A2 (n_1152));
AOI21_X1 i_1906 (.ZN (n_1384), .A (n_1376), .B1 (n_1382), .B2 (n_1383));
AND2_X1 i_1905 (.ZN (n_1383), .A1 (A[19]), .A2 (B[5]));
NOR2_X1 i_1904 (.ZN (n_1382), .A1 (n_1381), .A2 (n_1376));
AOI22_X1 i_1903 (.ZN (n_1381), .A1 (n_1377), .A2 (A[21]), .B1 (n_1378), .B2 (A[20]));
INV_X1 i_1902 (.ZN (n_1378), .A (n_340));
INV_X1 i_1901 (.ZN (n_1377), .A (n_424));
NOR3_X1 i_1900 (.ZN (n_1376), .A1 (n_1317), .A2 (n_1194), .A3 (n_340));
NAND2_X1 i_1899 (.ZN (n_1375), .A1 (B[7]), .A2 (A[18]));
XNOR2_X1 i_1898 (.ZN (n_1374), .A (n_1366), .B (n_1373));
OAI21_X1 i_1897 (.ZN (n_1373), .A (n_1369), .B1 (n_1371), .B2 (n_1372));
NAND2_X1 i_1896 (.ZN (n_1372), .A1 (A[2]), .A2 (B[23]));
NAND2_X1 i_1895 (.ZN (n_1371), .A1 (n_1369), .A2 (n_1370));
OAI22_X1 i_1894 (.ZN (n_1370), .A1 (n_1367), .A2 (n_422), .B1 (n_1368), .B2 (n_99));
NAND4_X1 i_1893 (.ZN (n_1369), .A1 (A[4]), .A2 (A[3]), .A3 (B[21]), .A4 (B[22]));
INV_X1 i_1892 (.ZN (n_1368), .A (B[22]));
INV_X1 i_1891 (.ZN (n_1367), .A (B[21]));
AOI22_X1 i_1890 (.ZN (n_1366), .A1 (n_1365), .A2 (n_1362), .B1 (n_1361), .B2 (n_1349));
OAI33_X1 i_1889 (.ZN (n_1365), .A1 (n_1364), .A2 (n_556), .A3 (n_1232), .B1 (n_458)
    , .B2 (n_592), .B3 (n_1363));
XNOR2_X1 i_1888 (.ZN (n_1364), .A (n_1363), .B (n_1230));
NAND2_X1 i_1887 (.ZN (n_1363), .A1 (A[9]), .A2 (B[15]));
XOR2_X1 i_1886 (.Z (n_1362), .A (n_1349), .B (n_1361));
OAI21_X1 i_1885 (.ZN (n_1361), .A (n_1358), .B1 (n_1360), .B2 (n_1164));
OR2_X1 i_1884 (.ZN (n_1360), .A1 (n_1357), .A2 (n_1359));
AOI22_X1 i_1883 (.ZN (n_1359), .A1 (A[14]), .A2 (B[10]), .B1 (A[15]), .B2 (B[9]));
INV_X1 i_1882 (.ZN (n_1358), .A (n_1357));
NOR2_X1 i_1881 (.ZN (n_1357), .A1 (n_1344), .A2 (n_1157));
OAI21_X1 i_1880 (.ZN (n_1349), .A (n_1345), .B1 (n_1348), .B2 (n_1343));
NAND2_X1 i_1879 (.ZN (n_1348), .A1 (n_1345), .A2 (n_1346));
OAI22_X1 i_1878 (.ZN (n_1346), .A1 (n_1339), .A2 (n_559), .B1 (n_229), .B2 (n_1235));
OR3_X1 i_1877 (.ZN (n_1345), .A1 (n_1341), .A2 (n_1339), .A3 (n_229));
NAND2_X1 i_1876 (.ZN (n_1344), .A1 (B[10]), .A2 (A[15]));
NAND2_X1 i_1875 (.ZN (n_1343), .A1 (A[12]), .A2 (B[12]));
NAND2_X1 i_1874 (.ZN (n_1341), .A1 (A[11]), .A2 (B[14]));
INV_X1 i_1873 (.ZN (n_1339), .A (A[10]));
AOI21_X1 i_1872 (.ZN (n_1338), .A (n_1330), .B1 (n_1332), .B2 (n_1334));
NOR2_X1 i_1871 (.ZN (n_1334), .A1 (n_1330), .A2 (n_1333));
AOI22_X1 i_1870 (.ZN (n_1333), .A1 (A[22]), .A2 (B[2]), .B1 (A[23]), .B2 (B[1]));
AOI21_X1 i_1869 (.ZN (n_1332), .A (n_1327), .B1 (n_1331), .B2 (n_949));
INV_X1 i_1868 (.ZN (n_1331), .A (n_1329));
NOR2_X1 i_1867 (.ZN (n_1330), .A1 (n_1328), .A2 (n_949));
NOR2_X1 i_1866 (.ZN (n_1329), .A1 (n_1328), .A2 (n_988));
NAND2_X1 i_1865 (.ZN (n_1328), .A1 (B[2]), .A2 (A[23]));
AOI22_X1 i_1864 (.ZN (n_1327), .A1 (A[21]), .A2 (B[2]), .B1 (B[0]), .B2 (A[23]));
XNOR2_X1 i_1863 (.ZN (n_1326), .A (n_1324), .B (n_1325));
AOI22_X1 i_1862 (.ZN (n_1325), .A1 (n_1190), .A2 (n_1154), .B1 (n_1153), .B2 (n_1147));
XNOR2_X1 i_1861 (.ZN (n_1324), .A (n_1321), .B (n_1323));
NOR2_X1 i_1860 (.ZN (n_1323), .A1 (n_1322), .A2 (n_1029));
INV_X1 i_1859 (.ZN (n_1322), .A (A[20]));
NOR2_X1 i_1858 (.ZN (n_1321), .A1 (n_1319), .A2 (n_1320));
AOI22_X1 i_1857 (.ZN (n_1320), .A1 (B[3]), .A2 (A[22]), .B1 (B[4]), .B2 (A[21]));
NOR3_X1 i_1856 (.ZN (n_1319), .A1 (n_1318), .A2 (n_1317), .A3 (n_424));
NAND2_X1 i_1855 (.ZN (n_1318), .A1 (B[4]), .A2 (A[22]));
INV_X1 i_1854 (.ZN (n_1317), .A (A[21]));
INV_X1 i_1853 (.ZN (n_1305), .A (A[16]));
OR3_X1 i_1852 (.ZN (n_1303), .A1 (n_1152), .A2 (n_1029), .A3 (n_1305));
OAI22_X1 i_1851 (.ZN (n_1302), .A1 (n_1305), .A2 (n_169), .B1 (n_1029), .B2 (n_1027));
NAND2_X1 i_1850 (.ZN (n_1301), .A1 (n_1303), .A2 (n_1302));
NAND2_X1 i_1849 (.ZN (n_1300), .A1 (A[15]), .A2 (B[7]));
OR2_X1 i_1848 (.ZN (n_1299), .A1 (n_954), .A2 (n_1194));
AOI22_X1 i_1847 (.ZN (n_1298), .A1 (A[20]), .A2 (B[2]), .B1 (A[19]), .B2 (B[3]));
INV_X1 i_1846 (.ZN (n_1297), .A (n_1298));
NAND2_X1 i_1845 (.ZN (n_1296), .A1 (n_1299), .A2 (n_1297));
NAND2_X1 i_1844 (.ZN (n_1295), .A1 (A[18]), .A2 (B[4]));
OAI21_X1 i_1843 (.ZN (n_1294), .A (n_1303), .B1 (n_1301), .B2 (n_1300));
OAI21_X1 i_1842 (.ZN (n_1293), .A (n_1299), .B1 (n_1296), .B2 (n_1295));
XOR2_X1 i_1841 (.Z (n_1292), .A (n_1294), .B (n_1293));
NOR2_X1 i_1840 (.ZN (n_1291), .A1 (n_1016), .A2 (n_1157));
AOI22_X1 i_1839 (.ZN (n_1290), .A1 (A[13]), .A2 (B[9]), .B1 (A[14]), .B2 (B[8]));
NOR2_X1 i_1838 (.ZN (n_1289), .A1 (n_1291), .A2 (n_1290));
OAI22_X1 i_1837 (.ZN (n_1266), .A1 (n_1016), .A2 (n_1157), .B1 (n_1173), .B2 (n_1290));
INV_X1 i_1836 (.ZN (n_1264), .A (n_1266));
AOI22_X1 i_1835 (.ZN (n_1263), .A1 (n_1294), .A2 (n_1293), .B1 (n_1292), .B2 (n_1266));
NAND2_X1 i_1834 (.ZN (n_1262), .A1 (A[2]), .A2 (B[21]));
NAND2_X1 i_1833 (.ZN (n_1261), .A1 (A[1]), .A2 (B[22]));
XNOR2_X1 i_1832 (.ZN (n_1260), .A (n_1262), .B (n_1261));
NAND2_X1 i_1831 (.ZN (n_1259), .A1 (A[0]), .A2 (B[23]));
OAI22_X1 i_1830 (.ZN (n_1239), .A1 (n_1262), .A2 (n_1261), .B1 (n_1260), .B2 (n_1259));
XNOR2_X1 i_1829 (.ZN (n_1236), .A (n_1263), .B (n_1239));
INV_X1 i_1828 (.ZN (n_1235), .A (A[11]));
INV_X1 i_1827 (.ZN (n_1232), .A (B[17]));
NAND2_X1 i_1826 (.ZN (n_1231), .A1 (A[7]), .A2 (B[15]));
NAND2_X1 i_1825 (.ZN (n_1230), .A1 (A[8]), .A2 (B[16]));
NOR2_X1 i_1824 (.ZN (n_1228), .A1 (n_1231), .A2 (n_1230));
AOI22_X1 i_1823 (.ZN (n_1227), .A1 (A[8]), .A2 (B[15]), .B1 (A[7]), .B2 (B[16]));
NOR2_X1 i_1822 (.ZN (n_1226), .A1 (n_1228), .A2 (n_1227));
NOR2_X1 i_1821 (.ZN (n_1225), .A1 (n_1232), .A2 (n_170));
AOI21_X1 i_1820 (.ZN (n_1222), .A (n_1228), .B1 (n_1226), .B2 (n_1225));
AOI22_X1 i_1819 (.ZN (n_1221), .A1 (A[10]), .A2 (B[13]), .B1 (A[11]), .B2 (B[12]));
OR3_X1 i_1818 (.ZN (n_1220), .A1 (n_1235), .A2 (n_229), .A3 (n_1060));
NAND2_X1 i_1817 (.ZN (n_1214), .A1 (A[9]), .A2 (B[14]));
AOI21_X1 i_1816 (.ZN (n_1213), .A (n_1221), .B1 (n_1220), .B2 (n_1214));
XNOR2_X1 i_1815 (.ZN (n_1212), .A (n_1222), .B (n_1213));
NAND2_X1 i_1814 (.ZN (n_1209), .A1 (A[4]), .A2 (B[18]));
NAND2_X1 i_1813 (.ZN (n_1205), .A1 (A[5]), .A2 (B[19]));
AOI22_X1 i_1812 (.ZN (n_1204), .A1 (A[5]), .A2 (B[18]), .B1 (A[4]), .B2 (B[19]));
INV_X1 i_1811 (.ZN (n_1203), .A (n_1204));
OAI21_X1 i_1810 (.ZN (n_1200), .A (n_1203), .B1 (n_1209), .B2 (n_1205));
NAND2_X1 i_1809 (.ZN (n_1199), .A1 (A[3]), .A2 (B[20]));
OAI22_X1 i_1808 (.ZN (n_1198), .A1 (n_1209), .A2 (n_1205), .B1 (n_1200), .B2 (n_1199));
XOR2_X1 i_1807 (.Z (n_1197), .A (n_1212), .B (n_1198));
INV_X1 i_1806 (.ZN (n_1196), .A (n_1197));
NAND2_X1 i_1805 (.ZN (n_1194), .A1 (A[20]), .A2 (B[3]));
NAND2_X1 i_1804 (.ZN (n_1193), .A1 (A[19]), .A2 (B[4]));
XNOR2_X1 i_1803 (.ZN (n_1192), .A (n_1194), .B (n_1193));
NAND2_X1 i_1802 (.ZN (n_1191), .A1 (A[18]), .A2 (B[5]));
OAI22_X1 i_1801 (.ZN (n_1190), .A1 (n_1194), .A2 (n_1193), .B1 (n_1192), .B2 (n_1191));
NAND2_X1 i_1800 (.ZN (n_1173), .A1 (A[12]), .A2 (B[10]));
NAND2_X1 i_1799 (.ZN (n_1164), .A1 (A[13]), .A2 (B[11]));
NOR2_X1 i_1798 (.ZN (n_1161), .A1 (n_1173), .A2 (n_1164));
INV_X1 i_1797 (.ZN (n_1160), .A (n_1161));
AOI22_X1 i_1796 (.ZN (n_1159), .A1 (A[12]), .A2 (B[11]), .B1 (A[13]), .B2 (B[10]));
NOR2_X1 i_1795 (.ZN (n_1158), .A1 (n_1161), .A2 (n_1159));
NAND2_X1 i_1794 (.ZN (n_1157), .A1 (A[14]), .A2 (B[9]));
AOI21_X1 i_1793 (.ZN (n_1154), .A (n_1159), .B1 (n_1160), .B2 (n_1157));
XOR2_X1 i_1792 (.Z (n_1153), .A (n_1190), .B (n_1154));
NAND2_X1 i_1791 (.ZN (n_1152), .A1 (A[17]), .A2 (B[6]));
NAND2_X1 i_1790 (.ZN (n_1151), .A1 (A[16]), .A2 (B[7]));
XNOR2_X1 i_1789 (.ZN (n_1150), .A (n_1152), .B (n_1151));
NAND2_X1 i_1788 (.ZN (n_1148), .A1 (A[15]), .A2 (B[8]));
OAI22_X1 i_1787 (.ZN (n_1147), .A1 (n_1152), .A2 (n_1151), .B1 (n_1150), .B2 (n_1148));
XOR2_X1 i_1786 (.Z (n_1146), .A (n_1153), .B (n_1147));
INV_X1 i_1785 (.ZN (n_1145), .A (n_1146));
AOI22_X1 i_1784 (.ZN (n_1144), .A1 (n_1197), .A2 (n_1146), .B1 (n_1196), .B2 (n_1145));
INV_X1 i_1783 (.ZN (n_1143), .A (n_837));
INV_X1 i_1782 (.ZN (n_1129), .A (n_953));
NAND2_X1 i_1781 (.ZN (n_1128), .A1 (B[5]), .A2 (A[13]));
NOR2_X1 i_1780 (.ZN (n_1122), .A1 (n_1011), .A2 (n_1128));
AOI22_X1 i_1779 (.ZN (n_1121), .A1 (B[5]), .A2 (A[14]), .B1 (B[6]), .B2 (A[13]));
NOR2_X1 i_1778 (.ZN (n_1120), .A1 (n_1122), .A2 (n_1121));
OAI22_X1 i_1777 (.ZN (n_1119), .A1 (n_1011), .A2 (n_1128), .B1 (n_1017), .B2 (n_1121));
AOI21_X1 i_1776 (.ZN (n_1118), .A (n_1143), .B1 (n_836), .B2 (n_838));
XOR2_X1 i_1775 (.Z (n_1117), .A (n_1119), .B (n_1118));
NAND2_X1 i_1774 (.ZN (n_1116), .A1 (B[8]), .A2 (A[11]));
XNOR2_X1 i_1773 (.ZN (n_1115), .A (n_1026), .B (n_1116));
NAND2_X1 i_1772 (.ZN (n_1114), .A1 (B[10]), .A2 (A[9]));
OAI22_X1 i_1771 (.ZN (n_1113), .A1 (n_1026), .A2 (n_1116), .B1 (n_1115), .B2 (n_1114));
NOR2_X1 i_1770 (.ZN (n_1112), .A1 (n_952), .A2 (n_1129));
XOR2_X1 i_1769 (.Z (n_1111), .A (n_951), .B (n_1112));
AOI22_X1 i_1768 (.ZN (n_1110), .A1 (n_1119), .A2 (n_1118), .B1 (n_1117), .B2 (n_1113));
INV_X1 i_1767 (.ZN (n_1104), .A (n_1110));
XOR2_X1 i_1766 (.Z (n_1103), .A (n_1111), .B (n_1104));
NAND2_X1 i_1765 (.ZN (n_1102), .A1 (B[4]), .A2 (A[17]));
NAND2_X1 i_1764 (.ZN (n_1101), .A1 (B[5]), .A2 (A[16]));
AND2_X1 i_1763 (.ZN (n_1100), .A1 (n_1102), .A2 (n_1101));
XOR2_X1 i_1762 (.Z (n_1099), .A (n_1102), .B (n_1101));
NAND2_X1 i_1761 (.ZN (n_1098), .A1 (B[6]), .A2 (A[15]));
XNOR2_X1 i_1760 (.ZN (n_1097), .A (n_1099), .B (n_1098));
AOI22_X1 i_1759 (.ZN (n_1096), .A1 (n_1111), .A2 (n_1104), .B1 (n_1103), .B2 (n_1097));
NAND2_X1 i_1758 (.ZN (n_1095), .A1 (B[7]), .A2 (A[14]));
XNOR2_X1 i_1757 (.ZN (n_1065), .A (n_1016), .B (n_1095));
NAND2_X1 i_1756 (.ZN (n_1064), .A1 (B[9]), .A2 (A[12]));
OAI22_X1 i_1755 (.ZN (n_1063), .A1 (n_1016), .A2 (n_1095), .B1 (n_1065), .B2 (n_1064));
OAI22_X1 i_1754 (.ZN (n_1062), .A1 (n_1102), .A2 (n_1101), .B1 (n_1100), .B2 (n_1098));
XOR2_X1 i_1753 (.Z (n_1061), .A (n_1063), .B (n_1062));
NAND2_X1 i_1752 (.ZN (n_1060), .A1 (B[12]), .A2 (A[10]));
AOI22_X1 i_1751 (.ZN (n_1059), .A1 (B[12]), .A2 (A[9]), .B1 (B[11]), .B2 (A[10]));
INV_X1 i_1750 (.ZN (n_1058), .A (n_1059));
OAI21_X1 i_1749 (.ZN (n_1057), .A (n_1058), .B1 (n_1021), .B2 (n_1060));
OAI22_X1 i_1748 (.ZN (n_1056), .A1 (n_1021), .A2 (n_1060), .B1 (n_1025), .B2 (n_1057));
XNOR2_X1 i_1747 (.ZN (n_1055), .A (n_1065), .B (n_1064));
XNOR2_X1 i_1746 (.ZN (n_1054), .A (n_1025), .B (n_1057));
NAND2_X1 i_1745 (.ZN (n_1053), .A1 (n_1055), .A2 (n_1054));
NOR2_X1 i_1744 (.ZN (n_1052), .A1 (n_1055), .A2 (n_1054));
NAND2_X1 i_1743 (.ZN (n_1051), .A1 (B[14]), .A2 (A[8]));
NOR2_X1 i_1742 (.ZN (n_1050), .A1 (n_1007), .A2 (n_1051));
AOI22_X1 i_1741 (.ZN (n_1049), .A1 (B[13]), .A2 (A[8]), .B1 (B[14]), .B2 (A[7]));
NOR2_X1 i_1740 (.ZN (n_1048), .A1 (n_1050), .A2 (n_1049));
NOR2_X1 i_1739 (.ZN (n_1036), .A1 (n_170), .A2 (n_560));
XOR2_X1 i_1738 (.Z (n_1035), .A (n_1048), .B (n_1036));
OAI21_X1 i_1737 (.ZN (n_1034), .A (n_1053), .B1 (n_1052), .B2 (n_1035));
XNOR2_X1 i_1736 (.ZN (n_1033), .A (n_1061), .B (n_1056));
XOR2_X1 i_1735 (.Z (n_1032), .A (n_1034), .B (n_1033));
AOI22_X1 i_1734 (.ZN (n_1031), .A1 (n_1034), .A2 (n_1033), .B1 (n_1096), .B2 (n_1032));
INV_X1 i_1733 (.ZN (n_1030), .A (n_1031));
INV_X1 i_1732 (.ZN (n_1029), .A (B[5]));
INV_X1 i_1731 (.ZN (n_1028), .A (A[18]));
INV_X1 i_1730 (.ZN (n_1027), .A (A[17]));
NAND2_X1 i_1729 (.ZN (n_1026), .A1 (B[9]), .A2 (A[10]));
NAND2_X1 i_1728 (.ZN (n_1025), .A1 (B[10]), .A2 (A[11]));
NOR2_X1 i_1727 (.ZN (n_1024), .A1 (n_1026), .A2 (n_1025));
AOI22_X1 i_1726 (.ZN (n_1023), .A1 (B[9]), .A2 (A[11]), .B1 (B[10]), .B2 (A[10]));
NOR2_X1 i_1725 (.ZN (n_1022), .A1 (n_1024), .A2 (n_1023));
NAND2_X1 i_1724 (.ZN (n_1021), .A1 (B[11]), .A2 (A[9]));
INV_X1 i_1723 (.ZN (n_1018), .A (n_1021));
NAND2_X1 i_1722 (.ZN (n_1017), .A1 (B[7]), .A2 (A[12]));
NAND2_X1 i_1721 (.ZN (n_1016), .A1 (B[8]), .A2 (A[13]));
NOR2_X1 i_1720 (.ZN (n_1015), .A1 (n_1017), .A2 (n_1016));
AOI22_X1 i_1719 (.ZN (n_1014), .A1 (B[8]), .A2 (A[12]), .B1 (B[7]), .B2 (A[13]));
NOR2_X1 i_1718 (.ZN (n_1013), .A1 (n_1015), .A2 (n_1014));
NAND2_X1 i_1717 (.ZN (n_1011), .A1 (B[6]), .A2 (A[14]));
INV_X1 i_1716 (.ZN (n_1009), .A (n_1011));
NAND2_X1 i_1715 (.ZN (n_1008), .A1 (B[12]), .A2 (A[8]));
NAND2_X1 i_1714 (.ZN (n_1007), .A1 (B[13]), .A2 (A[7]));
AOI21_X1 i_1713 (.ZN (n_1006), .A (n_1024), .B1 (n_1022), .B2 (n_1018));
AOI21_X1 i_1712 (.ZN (n_1005), .A (n_1015), .B1 (n_1013), .B2 (n_1009));
NOR2_X1 i_1711 (.ZN (n_1004), .A1 (n_1006), .A2 (n_1005));
XNOR2_X1 i_1710 (.ZN (n_1003), .A (n_1008), .B (n_1007));
NAND2_X1 i_1709 (.ZN (n_1002), .A1 (B[14]), .A2 (A[6]));
OAI22_X1 i_1708 (.ZN (n_1001), .A1 (n_1008), .A2 (n_1007), .B1 (n_1003), .B2 (n_1002));
AOI21_X1 i_1707 (.ZN (n_1000), .A (n_1004), .B1 (n_1006), .B2 (n_1005));
AOI21_X1 i_1706 (.ZN (n_999), .A (n_1004), .B1 (n_1001), .B2 (n_1000));
NOR3_X1 i_1705 (.ZN (n_998), .A1 (n_839), .A2 (n_340), .A3 (n_1027));
AOI22_X1 i_1704 (.ZN (n_996), .A1 (B[3]), .A2 (A[17]), .B1 (B[4]), .B2 (A[16]));
NOR2_X1 i_1703 (.ZN (n_995), .A1 (n_998), .A2 (n_996));
NOR2_X1 i_1702 (.ZN (n_994), .A1 (n_1029), .A2 (n_558));
NAND2_X1 i_1701 (.ZN (n_993), .A1 (B[1]), .A2 (A[20]));
NOR3_X1 i_1700 (.ZN (n_992), .A1 (n_28), .A2 (n_993), .A3 (n_853));
AOI22_X1 i_1699 (.ZN (n_991), .A1 (B[0]), .A2 (A[20]), .B1 (B[1]), .B2 (A[19]));
NOR2_X1 i_1698 (.ZN (n_990), .A1 (n_992), .A2 (n_991));
NOR2_X1 i_1697 (.ZN (n_989), .A1 (n_1028), .A2 (n_29));
NAND2_X1 i_1696 (.ZN (n_988), .A1 (B[0]), .A2 (A[21]));
AOI21_X1 i_1695 (.ZN (n_987), .A (n_998), .B1 (n_995), .B2 (n_994));
AOI21_X1 i_1694 (.ZN (n_986), .A (n_992), .B1 (n_990), .B2 (n_989));
NAND2_X1 i_1693 (.ZN (n_985), .A1 (n_987), .A2 (n_986));
INV_X1 i_1692 (.ZN (n_984), .A (n_985));
OAI22_X1 i_1691 (.ZN (n_978), .A1 (n_987), .A2 (n_986), .B1 (n_988), .B2 (n_984));
XNOR2_X1 i_1690 (.ZN (n_955), .A (n_999), .B (n_978));
NAND2_X1 i_1689 (.ZN (n_954), .A1 (B[2]), .A2 (A[19]));
NAND2_X1 i_1688 (.ZN (n_953), .A1 (n_993), .A2 (n_954));
NOR2_X1 i_1687 (.ZN (n_952), .A1 (n_993), .A2 (n_954));
NOR2_X1 i_1686 (.ZN (n_951), .A1 (n_1028), .A2 (n_424));
OAI21_X1 i_1685 (.ZN (n_950), .A (n_953), .B1 (n_952), .B2 (n_951));
NAND2_X1 i_1684 (.ZN (n_949), .A1 (B[1]), .A2 (A[22]));
NOR2_X1 i_1683 (.ZN (n_948), .A1 (n_988), .A2 (n_949));
AOI22_X1 i_1682 (.ZN (n_947), .A1 (B[0]), .A2 (A[22]), .B1 (B[1]), .B2 (A[21]));
OR2_X1 i_1681 (.ZN (n_946), .A1 (n_948), .A2 (n_947));
XOR2_X1 i_1680 (.Z (n_945), .A (n_950), .B (n_946));
XNOR2_X1 i_1679 (.ZN (n_944), .A (n_955), .B (n_945));
XOR2_X1 i_1678 (.Z (n_943), .A (n_1001), .B (n_1000));
OAI21_X1 i_1677 (.ZN (n_942), .A (n_985), .B1 (n_987), .B2 (n_986));
XOR2_X1 i_1676 (.Z (n_941), .A (n_988), .B (n_942));
XOR2_X1 i_1675 (.Z (n_940), .A (n_943), .B (n_941));
NAND2_X1 i_1674 (.ZN (n_939), .A1 (B[16]), .A2 (A[4]));
NAND2_X1 i_1673 (.ZN (n_938), .A1 (B[15]), .A2 (A[5]));
XOR2_X1 i_1672 (.Z (n_929), .A (n_939), .B (n_938));
INV_X1 i_1671 (.ZN (n_928), .A (n_929));
XNOR2_X1 i_1670 (.ZN (n_927), .A (n_1003), .B (n_1002));
NAND2_X1 i_1669 (.ZN (n_926), .A1 (B[17]), .A2 (A[3]));
XOR2_X1 i_1668 (.Z (n_925), .A (n_929), .B (n_926));
XOR2_X1 i_1667 (.Z (n_924), .A (n_927), .B (n_925));
NAND2_X1 i_1666 (.ZN (n_913), .A1 (B[18]), .A2 (A[1]));
NOR2_X1 i_1665 (.ZN (n_912), .A1 (n_855), .A2 (n_913));
AOI22_X1 i_1664 (.ZN (n_911), .A1 (B[18]), .A2 (A[2]), .B1 (B[19]), .B2 (A[1]));
NOR2_X1 i_1663 (.ZN (n_910), .A1 (n_912), .A2 (n_911));
NAND2_X1 i_1662 (.ZN (n_909), .A1 (n_857), .A2 (n_910));
OAI21_X1 i_1661 (.ZN (n_906), .A (n_909), .B1 (n_857), .B2 (n_910));
AOI22_X1 i_1660 (.ZN (n_905), .A1 (n_927), .A2 (n_925), .B1 (n_924), .B2 (n_906));
AOI22_X1 i_1659 (.ZN (n_904), .A1 (n_943), .A2 (n_941), .B1 (n_940), .B2 (n_905));
XOR2_X1 i_1658 (.Z (n_903), .A (n_944), .B (n_904));
INV_X1 i_1657 (.ZN (n_902), .A (n_897));
XOR2_X1 i_1656 (.Z (n_901), .A (n_899), .B (n_887));
XNOR2_X1 i_1655 (.ZN (n_899), .A (n_898), .B (n_888));
NOR2_X1 i_1654 (.ZN (n_898), .A1 (n_897), .A2 (n_896));
NOR3_X1 i_1653 (.ZN (n_897), .A1 (n_889), .A2 (n_422), .A3 (n_592));
AOI22_X1 i_1652 (.ZN (n_896), .A1 (B[16]), .A2 (A[5]), .B1 (B[17]), .B2 (A[4]));
NAND2_X1 i_1651 (.ZN (n_889), .A1 (A[5]), .A2 (B[17]));
NAND2_X1 i_1650 (.ZN (n_888), .A1 (B[18]), .A2 (A[3]));
XNOR2_X1 i_1649 (.ZN (n_887), .A (n_886), .B (n_855));
NOR2_X1 i_1648 (.ZN (n_886), .A1 (n_885), .A2 (n_884));
INV_X1 i_1647 (.ZN (n_885), .A (n_860));
AOI22_X1 i_1646 (.ZN (n_884), .A1 (B[20]), .A2 (A[1]), .B1 (B[21]), .B2 (A[0]));
NAND3_X1 i_1645 (.ZN (n_860), .A1 (n_857), .A2 (A[1]), .A3 (B[21]));
NOR2_X1 i_1644 (.ZN (n_857), .A1 (n_856), .A2 (n_31));
INV_X1 i_1643 (.ZN (n_856), .A (B[20]));
NAND2_X1 i_1642 (.ZN (n_855), .A1 (B[19]), .A2 (A[2]));
INV_X1 i_1641 (.ZN (n_853), .A (A[19]));
OAI22_X1 i_1640 (.ZN (n_852), .A1 (n_612), .A2 (n_616), .B1 (n_640), .B2 (n_645));
OAI22_X1 i_1639 (.ZN (n_851), .A1 (n_667), .A2 (n_668), .B1 (n_669), .B2 (n_670));
NAND2_X1 i_1638 (.ZN (n_850), .A1 (n_852), .A2 (n_851));
OAI21_X1 i_1637 (.ZN (n_849), .A (n_850), .B1 (n_852), .B2 (n_851));
NAND2_X1 i_1636 (.ZN (n_848), .A1 (B[0]), .A2 (A[18]));
OAI21_X1 i_1635 (.ZN (n_847), .A (n_850), .B1 (n_849), .B2 (n_848));
AOI21_X1 i_1634 (.ZN (n_846), .A (n_696), .B1 (n_731), .B2 (n_737));
NOR3_X1 i_1633 (.ZN (n_845), .A1 (n_257), .A2 (n_848), .A3 (n_853));
INV_X1 i_1632 (.ZN (n_844), .A (n_845));
AOI22_X1 i_1631 (.ZN (n_843), .A1 (B[0]), .A2 (A[19]), .B1 (B[1]), .B2 (A[18]));
NOR2_X1 i_1630 (.ZN (n_842), .A1 (n_845), .A2 (n_843));
XNOR2_X1 i_1629 (.ZN (n_841), .A (n_846), .B (n_842));
XOR2_X1 i_1628 (.Z (n_840), .A (n_847), .B (n_841));
NAND2_X1 i_1627 (.ZN (n_839), .A1 (B[3]), .A2 (A[16]));
OR2_X1 i_1626 (.ZN (n_838), .A1 (n_695), .A2 (n_839));
NAND2_X1 i_1625 (.ZN (n_837), .A1 (n_695), .A2 (n_839));
NAND2_X1 i_1624 (.ZN (n_836), .A1 (B[4]), .A2 (A[15]));
NAND2_X1 i_1623 (.ZN (n_835), .A1 (n_838), .A2 (n_837));
XOR2_X1 i_1622 (.Z (n_834), .A (n_836), .B (n_835));
XNOR2_X1 i_1621 (.ZN (n_833), .A (n_840), .B (n_834));
OAI21_X1 i_1620 (.ZN (n_832), .A (n_830), .B1 (n_802), .B2 (n_831));
OAI21_X1 i_1619 (.ZN (n_831), .A (n_830), .B1 (n_829), .B2 (n_817));
NAND2_X1 i_1618 (.ZN (n_830), .A1 (n_817), .A2 (n_829));
OAI22_X1 i_1617 (.ZN (n_829), .A1 (n_666), .A2 (n_671), .B1 (n_664), .B2 (n_665));
XNOR2_X1 i_1616 (.ZN (n_817), .A (n_693), .B (n_761));
AOI21_X1 i_1615 (.ZN (n_802), .A (n_776), .B1 (n_777), .B2 (n_784));
INV_X1 i_1614 (.ZN (n_784), .A (n_783));
AOI22_X1 i_1613 (.ZN (n_783), .A1 (n_781), .A2 (n_782), .B1 (n_779), .B2 (n_780));
XOR2_X1 i_1612 (.Z (n_782), .A (n_676), .B (n_677));
XOR2_X1 i_1611 (.Z (n_781), .A (n_779), .B (n_780));
XOR2_X1 i_1610 (.Z (n_780), .A (n_682), .B (n_683));
XOR2_X1 i_1609 (.Z (n_779), .A (n_661), .B (n_778));
NOR2_X1 i_1608 (.ZN (n_778), .A1 (n_663), .A2 (n_647));
AOI21_X1 i_1607 (.ZN (n_777), .A (n_776), .B1 (n_774), .B2 (n_775));
NOR2_X1 i_1606 (.ZN (n_776), .A1 (n_774), .A2 (n_775));
XNOR2_X1 i_1605 (.ZN (n_775), .A (n_686), .B (n_692));
AOI21_X1 i_1604 (.ZN (n_774), .A (n_771), .B1 (n_772), .B2 (n_773));
XOR2_X1 i_1603 (.Z (n_773), .A (n_591), .B (n_593));
AOI21_X1 i_1602 (.ZN (n_772), .A (n_771), .B1 (n_770), .B2 (n_763));
NOR2_X1 i_1601 (.ZN (n_771), .A1 (n_763), .A2 (n_770));
XOR2_X1 i_1600 (.Z (n_770), .A (n_769), .B (n_601));
NOR2_X1 i_1599 (.ZN (n_769), .A1 (n_602), .A2 (n_600));
XNOR2_X1 i_1598 (.ZN (n_763), .A (n_762), .B (n_691));
NOR2_X1 i_1597 (.ZN (n_762), .A1 (n_687), .A2 (n_690));
XOR2_X1 i_1596 (.Z (n_761), .A (n_760), .B (n_750));
XNOR2_X1 i_1595 (.ZN (n_760), .A (n_731), .B (n_737));
OAI22_X1 i_1594 (.ZN (n_750), .A1 (n_608), .A2 (n_609), .B1 (n_583), .B2 (n_607));
NOR2_X1 i_1593 (.ZN (n_737), .A1 (n_424), .A2 (n_558));
NOR2_X1 i_1592 (.ZN (n_731), .A1 (n_696), .A2 (n_726));
AOI22_X1 i_1591 (.ZN (n_726), .A1 (A[16]), .A2 (B[2]), .B1 (A[17]), .B2 (B[1]));
NOR2_X1 i_1590 (.ZN (n_696), .A1 (n_612), .A2 (n_695));
NAND2_X1 i_1589 (.ZN (n_695), .A1 (B[2]), .A2 (A[17]));
INV_X1 i_1588 (.ZN (n_694), .A (n_693));
OAI21_X1 i_1587 (.ZN (n_693), .A (n_685), .B1 (n_686), .B2 (n_692));
OAI21_X1 i_1586 (.ZN (n_692), .A (n_689), .B1 (n_690), .B2 (n_691));
AND2_X1 i_1585 (.ZN (n_691), .A1 (A[6]), .A2 (B[10]));
NOR3_X1 i_1584 (.ZN (n_690), .A1 (n_567), .A2 (n_426), .A3 (n_458));
INV_X1 i_1583 (.ZN (n_689), .A (n_687));
AOI22_X1 i_1582 (.ZN (n_687), .A1 (A[7]), .A2 (B[9]), .B1 (A[8]), .B2 (B[8]));
OAI21_X1 i_1581 (.ZN (n_686), .A (n_685), .B1 (n_678), .B2 (n_684));
NAND2_X1 i_1580 (.ZN (n_685), .A1 (n_678), .A2 (n_684));
OAI21_X1 i_1579 (.ZN (n_684), .A (n_680), .B1 (n_682), .B2 (n_683));
OR2_X1 i_1578 (.ZN (n_683), .A1 (n_340), .A2 (n_258));
OR2_X1 i_1577 (.ZN (n_682), .A1 (n_679), .A2 (n_681));
AOI22_X1 i_1576 (.ZN (n_681), .A1 (A[13]), .A2 (B[3]), .B1 (A[14]), .B2 (B[2]));
INV_X1 i_1575 (.ZN (n_680), .A (n_679));
NOR2_X1 i_1574 (.ZN (n_679), .A1 (n_613), .A2 (n_667));
OAI22_X1 i_1573 (.ZN (n_678), .A1 (n_676), .A2 (n_677), .B1 (n_675), .B2 (n_561));
NAND2_X1 i_1572 (.ZN (n_677), .A1 (A[9]), .A2 (B[7]));
XNOR2_X1 i_1571 (.ZN (n_676), .A (n_675), .B (n_561));
NAND2_X1 i_1570 (.ZN (n_675), .A1 (A[10]), .A2 (B[6]));
XNOR2_X1 i_1569 (.ZN (n_671), .A (n_669), .B (n_670));
NAND2_X1 i_1568 (.ZN (n_670), .A1 (A[12]), .A2 (B[5]));
XNOR2_X1 i_1567 (.ZN (n_669), .A (n_667), .B (n_668));
NAND2_X1 i_1566 (.ZN (n_668), .A1 (B[4]), .A2 (A[13]));
NAND2_X1 i_1565 (.ZN (n_667), .A1 (B[3]), .A2 (A[14]));
XNOR2_X1 i_1564 (.ZN (n_666), .A (n_664), .B (n_665));
XNOR2_X1 i_1563 (.ZN (n_665), .A (n_640), .B (n_645));
OAI21_X1 i_1562 (.ZN (n_664), .A (n_660), .B1 (n_661), .B2 (n_663));
NOR2_X1 i_1561 (.ZN (n_663), .A1 (n_612), .A2 (n_662));
INV_X1 i_1560 (.ZN (n_662), .A (n_488));
OAI22_X1 i_1559 (.ZN (n_661), .A1 (n_614), .A2 (n_615), .B1 (n_613), .B2 (n_469));
INV_X1 i_1558 (.ZN (n_660), .A (n_647));
AOI22_X1 i_1557 (.ZN (n_647), .A1 (B[0]), .A2 (A[16]), .B1 (A[15]), .B2 (B[1]));
NAND2_X1 i_1556 (.ZN (n_645), .A1 (A[15]), .A2 (B[2]));
XNOR2_X1 i_1555 (.ZN (n_640), .A (n_612), .B (n_616));
NAND2_X1 i_1554 (.ZN (n_616), .A1 (B[0]), .A2 (A[17]));
NAND2_X1 i_1553 (.ZN (n_615), .A1 (A[12]), .A2 (B[3]));
XNOR2_X1 i_1552 (.ZN (n_614), .A (n_613), .B (n_469));
NAND2_X1 i_1551 (.ZN (n_613), .A1 (A[13]), .A2 (B[2]));
NAND2_X1 i_1550 (.ZN (n_612), .A1 (A[16]), .A2 (B[1]));
XOR2_X1 i_1549 (.Z (n_611), .A (n_606), .B (n_610));
XNOR2_X1 i_1548 (.ZN (n_610), .A (n_608), .B (n_609));
NAND2_X1 i_1547 (.ZN (n_609), .A1 (B[17]), .A2 (A[0]));
XNOR2_X1 i_1546 (.ZN (n_608), .A (n_583), .B (n_607));
NAND2_X1 i_1545 (.ZN (n_607), .A1 (B[16]), .A2 (A[1]));
XOR2_X1 i_1544 (.Z (n_606), .A (n_582), .B (n_605));
XNOR2_X1 i_1543 (.ZN (n_605), .A (n_598), .B (n_604));
OAI21_X1 i_1542 (.ZN (n_604), .A (n_603), .B1 (n_600), .B2 (n_601));
INV_X1 i_1541 (.ZN (n_603), .A (n_602));
NOR2_X1 i_1540 (.ZN (n_602), .A1 (n_599), .A2 (n_535));
NAND2_X1 i_1539 (.ZN (n_601), .A1 (B[13]), .A2 (A[3]));
AOI22_X1 i_1538 (.ZN (n_600), .A1 (B[12]), .A2 (A[4]), .B1 (B[11]), .B2 (A[5]));
NAND2_X1 i_1537 (.ZN (n_599), .A1 (B[12]), .A2 (A[5]));
AOI21_X1 i_1536 (.ZN (n_598), .A (n_589), .B1 (n_591), .B2 (n_593));
NOR2_X1 i_1535 (.ZN (n_593), .A1 (n_592), .A2 (n_31));
INV_X1 i_1534 (.ZN (n_592), .A (B[16]));
NOR2_X1 i_1533 (.ZN (n_591), .A1 (n_589), .A2 (n_590));
AOI22_X1 i_1532 (.ZN (n_590), .A1 (B[15]), .A2 (A[1]), .B1 (B[14]), .B2 (A[2]));
NOR2_X1 i_1531 (.ZN (n_589), .A1 (n_583), .A2 (n_515));
NAND2_X1 i_1530 (.ZN (n_583), .A1 (B[15]), .A2 (A[2]));
AOI21_X1 i_1529 (.ZN (n_582), .A (n_575), .B1 (n_576), .B2 (n_581));
AOI21_X1 i_1528 (.ZN (n_581), .A (n_578), .B1 (n_579), .B2 (n_580));
NAND3_X1 i_1527 (.ZN (n_580), .A1 (n_577), .A2 (B[12]), .A3 (A[3]));
NAND2_X1 i_1526 (.ZN (n_579), .A1 (B[10]), .A2 (A[5]));
AOI21_X1 i_1525 (.ZN (n_578), .A (n_577), .B1 (B[12]), .B2 (A[3]));
INV_X1 i_1524 (.ZN (n_577), .A (n_535));
AOI21_X1 i_1523 (.ZN (n_576), .A (n_575), .B1 (n_572), .B2 (n_574));
NOR2_X1 i_1522 (.ZN (n_575), .A1 (n_572), .A2 (n_574));
OAI21_X1 i_1521 (.ZN (n_574), .A (n_568), .B1 (n_570), .B2 (n_573));
INV_X1 i_1520 (.ZN (n_573), .A (n_569));
AOI21_X1 i_1519 (.ZN (n_572), .A (n_562), .B1 (n_565), .B2 (n_566));
INV_X1 i_1518 (.ZN (n_571), .A (n_570));
NOR2_X1 i_1517 (.ZN (n_570), .A1 (n_567), .A2 (n_544));
NAND2_X1 i_1516 (.ZN (n_569), .A1 (B[9]), .A2 (A[6]));
NAND2_X1 i_1515 (.ZN (n_568), .A1 (n_567), .A2 (n_544));
NAND2_X1 i_1514 (.ZN (n_567), .A1 (B[8]), .A2 (A[7]));
NOR2_X1 i_1513 (.ZN (n_566), .A1 (n_169), .A2 (n_339));
NOR2_X1 i_1512 (.ZN (n_565), .A1 (n_562), .A2 (n_564));
AOI22_X1 i_1511 (.ZN (n_564), .A1 (B[5]), .A2 (A[10]), .B1 (B[4]), .B2 (A[11]));
NOR2_X1 i_1510 (.ZN (n_562), .A1 (n_561), .A2 (n_494));
NAND2_X1 i_1509 (.ZN (n_561), .A1 (B[5]), .A2 (A[11]));
INV_X1 i_1508 (.ZN (n_560), .A (B[15]));
INV_X1 i_1507 (.ZN (n_559), .A (B[14]));
INV_X1 i_1506 (.ZN (n_558), .A (A[15]));
INV_X1 i_1505 (.ZN (n_557), .A (A[14]));
INV_X1 i_1504 (.ZN (n_556), .A (A[7]));
INV_X1 i_1503 (.ZN (n_555), .A (n_287));
NAND2_X1 i_1502 (.ZN (n_544), .A1 (B[7]), .A2 (A[8]));
NOR3_X1 i_1501 (.ZN (n_543), .A1 (n_169), .A2 (n_544), .A3 (n_556));
AOI22_X1 i_1500 (.ZN (n_542), .A1 (B[7]), .A2 (A[7]), .B1 (B[6]), .B2 (A[8]));
NOR2_X1 i_1499 (.ZN (n_541), .A1 (n_543), .A2 (n_542));
NOR2_X1 i_1498 (.ZN (n_540), .A1 (n_170), .A2 (n_425));
AOI22_X1 i_1497 (.ZN (n_537), .A1 (B[11]), .A2 (A[3]), .B1 (B[10]), .B2 (A[4]));
INV_X1 i_1496 (.ZN (n_536), .A (n_537));
NAND2_X1 i_1495 (.ZN (n_535), .A1 (B[11]), .A2 (A[4]));
NOR2_X1 i_1494 (.ZN (n_534), .A1 (n_284), .A2 (n_535));
AOI21_X1 i_1493 (.ZN (n_533), .A (n_543), .B1 (n_541), .B2 (n_540));
OAI21_X1 i_1492 (.ZN (n_532), .A (n_536), .B1 (n_555), .B2 (n_534));
NAND2_X1 i_1491 (.ZN (n_531), .A1 (n_533), .A2 (n_532));
INV_X1 i_1490 (.ZN (n_530), .A (n_531));
OAI21_X1 i_1489 (.ZN (n_524), .A (n_531), .B1 (n_533), .B2 (n_532));
AOI22_X1 i_1488 (.ZN (n_523), .A1 (B[12]), .A2 (A[2]), .B1 (B[13]), .B2 (A[1]));
INV_X1 i_1487 (.ZN (n_522), .A (n_523));
NAND2_X1 i_1486 (.ZN (n_521), .A1 (B[13]), .A2 (A[2]));
NOR2_X1 i_1485 (.ZN (n_520), .A1 (n_204), .A2 (n_521));
NOR2_X1 i_1484 (.ZN (n_517), .A1 (n_559), .A2 (n_31));
OAI21_X1 i_1483 (.ZN (n_516), .A (n_522), .B1 (n_520), .B2 (n_517));
NAND2_X1 i_1482 (.ZN (n_515), .A1 (B[14]), .A2 (A[1]));
XNOR2_X1 i_1481 (.ZN (n_502), .A (n_521), .B (n_515));
OAI33_X1 i_1480 (.ZN (n_501), .A1 (n_560), .A2 (n_31), .A3 (n_502), .B1 (n_33), .B2 (n_229), .B3 (n_515));
OAI22_X1 i_1479 (.ZN (n_498), .A1 (n_533), .A2 (n_532), .B1 (n_530), .B2 (n_516));
NAND2_X1 i_1478 (.ZN (n_496), .A1 (n_501), .A2 (n_498));
OAI21_X1 i_1477 (.ZN (n_495), .A (n_496), .B1 (n_501), .B2 (n_498));
NAND2_X1 i_1476 (.ZN (n_494), .A1 (B[4]), .A2 (A[10]));
XNOR2_X1 i_1475 (.ZN (n_492), .A (n_311), .B (n_494));
NAND2_X1 i_1474 (.ZN (n_489), .A1 (B[5]), .A2 (A[9]));
NOR2_X1 i_1473 (.ZN (n_488), .A1 (n_558), .A2 (n_28));
OAI22_X1 i_1472 (.ZN (n_487), .A1 (n_311), .A2 (n_494), .B1 (n_492), .B2 (n_489));
XOR2_X1 i_1471 (.Z (n_470), .A (n_488), .B (n_487));
NAND2_X1 i_1470 (.ZN (n_469), .A1 (B[1]), .A2 (A[14]));
OR3_X1 i_1469 (.ZN (n_468), .A1 (n_28), .A2 (n_469), .A3 (n_256));
OAI22_X1 i_1468 (.ZN (n_467), .A1 (n_557), .A2 (n_28), .B1 (n_256), .B2 (n_257));
NAND2_X1 i_1467 (.ZN (n_466), .A1 (n_468), .A2 (n_467));
NAND2_X1 i_1466 (.ZN (n_465), .A1 (B[2]), .A2 (A[12]));
OAI21_X1 i_1465 (.ZN (n_462), .A (n_468), .B1 (n_466), .B2 (n_465));
AOI22_X1 i_1464 (.ZN (n_461), .A1 (n_488), .A2 (n_487), .B1 (n_470), .B2 (n_462));
OAI21_X1 i_1463 (.ZN (n_460), .A (n_496), .B1 (n_495), .B2 (n_461));
INV_X1 i_1462 (.ZN (n_459), .A (n_460));
INV_X1 i_1461 (.ZN (n_458), .A (A[8]));
INV_X1 i_1460 (.ZN (n_457), .A (n_338));
NAND2_X1 i_1459 (.ZN (n_455), .A1 (B[2]), .A2 (A[7]));
XNOR2_X1 i_1458 (.ZN (n_454), .A (n_420), .B (n_455));
OAI33_X1 i_1457 (.ZN (n_453), .A1 (n_424), .A2 (n_170), .A3 (n_454), .B1 (n_458), .B2 (n_257), .B3 (n_455));
XOR2_X1 i_1456 (.Z (n_446), .A (n_457), .B (n_453));
NOR2_X1 i_1455 (.ZN (n_445), .A1 (n_257), .A2 (n_339));
AOI22_X1 i_1454 (.ZN (n_444), .A1 (n_457), .A2 (n_453), .B1 (n_446), .B2 (n_445));
XNOR2_X1 i_1453 (.ZN (n_442), .A (n_333), .B (n_332));
NOR2_X1 i_1452 (.ZN (n_441), .A1 (n_444), .A2 (n_442));
AOI21_X1 i_1451 (.ZN (n_439), .A (n_441), .B1 (n_444), .B2 (n_442));
NAND2_X1 i_1450 (.ZN (n_438), .A1 (n_327), .A2 (n_330));
XOR2_X1 i_1449 (.Z (n_437), .A (n_328), .B (n_438));
AOI21_X1 i_1448 (.ZN (n_427), .A (n_441), .B1 (n_439), .B2 (n_437));
INV_X1 i_1447 (.ZN (n_426), .A (B[9]));
INV_X1 i_1446 (.ZN (n_425), .A (B[8]));
INV_X1 i_1445 (.ZN (n_424), .A (B[3]));
INV_X1 i_1444 (.ZN (n_423), .A (A[5]));
INV_X1 i_1443 (.ZN (n_422), .A (A[4]));
NAND2_X1 i_1442 (.ZN (n_421), .A1 (B[0]), .A2 (A[7]));
NAND2_X1 i_1441 (.ZN (n_420), .A1 (B[1]), .A2 (A[8]));
NOR2_X1 i_1440 (.ZN (n_419), .A1 (n_421), .A2 (n_420));
AOI22_X1 i_1439 (.ZN (n_418), .A1 (B[0]), .A2 (A[8]), .B1 (B[1]), .B2 (A[7]));
NOR2_X1 i_1438 (.ZN (n_417), .A1 (n_419), .A2 (n_418));
NOR2_X1 i_1437 (.ZN (n_416), .A1 (n_29), .A2 (n_170));
OR2_X1 i_1436 (.ZN (n_400), .A1 (n_28), .A2 (n_339));
AOI21_X1 i_1435 (.ZN (n_399), .A (n_419), .B1 (n_417), .B2 (n_416));
NOR2_X1 i_1434 (.ZN (n_398), .A1 (n_400), .A2 (n_399));
AOI21_X1 i_1433 (.ZN (n_397), .A (n_398), .B1 (n_400), .B2 (n_399));
NAND2_X1 i_1432 (.ZN (n_396), .A1 (B[4]), .A2 (A[5]));
OR3_X1 i_1431 (.ZN (n_395), .A1 (n_424), .A2 (n_396), .A3 (n_422));
OAI22_X1 i_1430 (.ZN (n_394), .A1 (n_424), .A2 (n_423), .B1 (n_422), .B2 (n_340));
NAND2_X1 i_1429 (.ZN (n_393), .A1 (n_395), .A2 (n_394));
NAND2_X1 i_1428 (.ZN (n_392), .A1 (B[5]), .A2 (A[3]));
OAI21_X1 i_1427 (.ZN (n_391), .A (n_395), .B1 (n_393), .B2 (n_392));
AOI21_X1 i_1426 (.ZN (n_390), .A (n_398), .B1 (n_397), .B2 (n_391));
NAND2_X1 i_1425 (.ZN (n_389), .A1 (B[5]), .A2 (A[4]));
XNOR2_X1 i_1424 (.ZN (n_388), .A (n_396), .B (n_389));
NAND2_X1 i_1423 (.ZN (n_387), .A1 (B[6]), .A2 (A[3]));
NAND2_X1 i_1422 (.ZN (n_386), .A1 (B[7]), .A2 (A[1]));
NAND2_X1 i_1421 (.ZN (n_385), .A1 (B[8]), .A2 (A[2]));
NOR2_X1 i_1420 (.ZN (n_384), .A1 (n_386), .A2 (n_385));
AOI22_X1 i_1419 (.ZN (n_382), .A1 (B[8]), .A2 (A[1]), .B1 (B[7]), .B2 (A[2]));
NOR2_X1 i_1418 (.ZN (n_381), .A1 (n_384), .A2 (n_382));
NOR2_X1 i_1417 (.ZN (n_380), .A1 (n_426), .A2 (n_31));
AOI21_X1 i_1416 (.ZN (n_379), .A (n_384), .B1 (n_381), .B2 (n_380));
OAI22_X1 i_1415 (.ZN (n_378), .A1 (n_396), .A2 (n_389), .B1 (n_388), .B2 (n_387));
INV_X1 i_1414 (.ZN (n_377), .A (n_378));
XNOR2_X1 i_1413 (.ZN (n_376), .A (n_379), .B (n_377));
OAI22_X1 i_1412 (.ZN (n_375), .A1 (n_379), .A2 (n_377), .B1 (n_390), .B2 (n_376));
NAND2_X1 i_1411 (.ZN (n_374), .A1 (B[9]), .A2 (A[1]));
NOR2_X1 i_1410 (.ZN (n_373), .A1 (n_208), .A2 (n_374));
AOI22_X1 i_1409 (.ZN (n_372), .A1 (B[9]), .A2 (A[2]), .B1 (B[10]), .B2 (A[1]));
NOR2_X1 i_1408 (.ZN (n_371), .A1 (n_373), .A2 (n_372));
NAND2_X1 i_1407 (.ZN (n_370), .A1 (B[6]), .A2 (A[4]));
NOR2_X1 i_1406 (.ZN (n_369), .A1 (n_175), .A2 (n_370));
AOI22_X1 i_1405 (.ZN (n_368), .A1 (B[6]), .A2 (A[5]), .B1 (B[7]), .B2 (A[4]));
NOR2_X1 i_1404 (.ZN (n_359), .A1 (n_369), .A2 (n_368));
NOR2_X1 i_1403 (.ZN (n_358), .A1 (n_425), .A2 (n_99));
XNOR2_X1 i_1402 (.ZN (n_357), .A (n_198), .B (n_371));
XOR2_X1 i_1401 (.Z (n_356), .A (n_359), .B (n_358));
XOR2_X1 i_1400 (.Z (n_355), .A (n_357), .B (n_356));
AOI22_X1 i_1399 (.ZN (n_354), .A1 (n_357), .A2 (n_356), .B1 (n_375), .B2 (n_355));
INV_X1 i_1398 (.ZN (n_340), .A (B[4]));
INV_X1 i_1397 (.ZN (n_339), .A (A[9]));
NAND2_X1 i_1396 (.ZN (n_338), .A1 (B[0]), .A2 (A[10]));
NOR2_X1 i_1395 (.ZN (n_335), .A1 (n_260), .A2 (n_338));
AOI22_X1 i_1394 (.ZN (n_334), .A1 (B[1]), .A2 (A[10]), .B1 (B[0]), .B2 (A[11]));
NOR2_X1 i_1393 (.ZN (n_333), .A1 (n_335), .A2 (n_334));
NOR2_X1 i_1392 (.ZN (n_332), .A1 (n_339), .A2 (n_29));
NAND2_X1 i_1391 (.ZN (n_331), .A1 (B[3]), .A2 (A[8]));
NAND2_X1 i_1390 (.ZN (n_330), .A1 (n_272), .A2 (n_331));
NAND2_X1 i_1389 (.ZN (n_328), .A1 (B[5]), .A2 (A[6]));
OR2_X1 i_1388 (.ZN (n_327), .A1 (n_272), .A2 (n_331));
AOI21_X1 i_1387 (.ZN (n_326), .A (n_335), .B1 (n_333), .B2 (n_332));
NAND2_X1 i_1386 (.ZN (n_325), .A1 (n_328), .A2 (n_327));
NAND2_X1 i_1385 (.ZN (n_324), .A1 (n_330), .A2 (n_325));
NOR2_X1 i_1384 (.ZN (n_323), .A1 (n_326), .A2 (n_324));
AOI21_X1 i_1383 (.ZN (n_321), .A (n_323), .B1 (n_326), .B2 (n_324));
NAND2_X1 i_1382 (.ZN (n_320), .A1 (n_265), .A2 (n_259));
XOR2_X1 i_1381 (.Z (n_319), .A (n_264), .B (n_320));
AOI21_X1 i_1380 (.ZN (n_314), .A (n_323), .B1 (n_269), .B2 (n_321));
NOR2_X1 i_1379 (.ZN (n_313), .A1 (n_319), .A2 (n_314));
AOI21_X1 i_1378 (.ZN (n_312), .A (n_313), .B1 (n_319), .B2 (n_314));
NAND2_X1 i_1377 (.ZN (n_311), .A1 (B[3]), .A2 (A[11]));
NOR2_X1 i_1376 (.ZN (n_309), .A1 (n_261), .A2 (n_311));
AOI22_X1 i_1375 (.ZN (n_308), .A1 (B[3]), .A2 (A[10]), .B1 (B[2]), .B2 (A[11]));
NOR2_X1 i_1374 (.ZN (n_307), .A1 (n_309), .A2 (n_308));
NOR2_X1 i_1373 (.ZN (n_306), .A1 (n_340), .A2 (n_339));
XOR2_X1 i_1372 (.Z (n_305), .A (n_307), .B (n_306));
AOI21_X1 i_1371 (.ZN (n_304), .A (n_313), .B1 (n_312), .B2 (n_305));
NAND2_X1 i_1370 (.ZN (n_287), .A1 (B[9]), .A2 (A[5]));
NOR2_X1 i_1369 (.ZN (n_286), .A1 (n_176), .A2 (n_287));
AOI22_X1 i_1368 (.ZN (n_285), .A1 (B[8]), .A2 (A[5]), .B1 (B[9]), .B2 (A[4]));
NAND2_X1 i_1367 (.ZN (n_284), .A1 (B[10]), .A2 (A[3]));
NAND3_X1 i_1366 (.ZN (n_283), .A1 (A[7]), .A2 (n_171), .A3 (B[7]));
INV_X1 i_1365 (.ZN (n_282), .A (n_283));
AOI22_X1 i_1364 (.ZN (n_281), .A1 (B[6]), .A2 (A[7]), .B1 (B[7]), .B2 (A[6]));
NOR2_X1 i_1363 (.ZN (n_280), .A1 (n_286), .A2 (n_285));
XOR2_X1 i_1362 (.Z (n_279), .A (n_284), .B (n_280));
NOR2_X1 i_1361 (.ZN (n_278), .A1 (n_282), .A2 (n_281));
XOR2_X1 i_1360 (.Z (n_277), .A (n_270), .B (n_278));
XOR2_X1 i_1359 (.Z (n_276), .A (n_279), .B (n_277));
XNOR2_X1 i_1358 (.ZN (n_275), .A (n_228), .B (n_230));
AOI22_X1 i_1357 (.ZN (n_274), .A1 (n_279), .A2 (n_277), .B1 (n_276), .B2 (n_275));
XNOR2_X1 i_1356 (.ZN (n_273), .A (n_304), .B (n_274));
NAND2_X1 i_1355 (.ZN (n_272), .A1 (B[4]), .A2 (A[7]));
NAND2_X1 i_1354 (.ZN (n_270), .A1 (B[5]), .A2 (A[8]));
NOR2_X1 i_1353 (.ZN (n_269), .A1 (n_258), .A2 (n_28));
XNOR2_X1 i_1352 (.ZN (n_268), .A (n_246), .B (n_267));
OAI21_X1 i_1351 (.ZN (n_267), .A (n_259), .B1 (n_264), .B2 (n_266));
INV_X1 i_1350 (.ZN (n_266), .A (n_265));
OR4_X1 i_1349 (.ZN (n_265), .A1 (n_256), .A2 (n_258), .A3 (n_257), .A4 (n_28));
OAI22_X1 i_1348 (.ZN (n_264), .A1 (n_262), .A2 (n_263), .B1 (n_260), .B2 (n_261));
NAND2_X1 i_1347 (.ZN (n_263), .A1 (B[3]), .A2 (A[9]));
XNOR2_X1 i_1346 (.ZN (n_262), .A (n_260), .B (n_261));
NAND2_X1 i_1345 (.ZN (n_261), .A1 (B[2]), .A2 (A[10]));
NAND2_X1 i_1344 (.ZN (n_260), .A1 (B[1]), .A2 (A[11]));
OAI22_X1 i_1343 (.ZN (n_259), .A1 (n_258), .A2 (n_257), .B1 (n_256), .B2 (n_28));
INV_X1 i_1342 (.ZN (n_258), .A (A[12]));
INV_X1 i_1341 (.ZN (n_257), .A (B[1]));
INV_X1 i_1340 (.ZN (n_256), .A (A[13]));
XNOR2_X1 i_1339 (.ZN (n_246), .A (n_222), .B (n_245));
AOI21_X1 i_1338 (.ZN (n_245), .A (n_227), .B1 (n_228), .B2 (n_230));
NOR2_X1 i_1337 (.ZN (n_230), .A1 (n_229), .A2 (n_31));
INV_X1 i_1336 (.ZN (n_229), .A (B[13]));
AOI21_X1 i_1335 (.ZN (n_228), .A (n_227), .B1 (n_204), .B2 (n_226));
NOR2_X1 i_1334 (.ZN (n_227), .A1 (n_204), .A2 (n_226));
NAND2_X1 i_1333 (.ZN (n_226), .A1 (B[11]), .A2 (A[2]));
OAI21_X1 i_1332 (.ZN (n_222), .A (n_188), .B1 (n_189), .B2 (n_212));
AOI21_X1 i_1331 (.ZN (n_212), .A (n_205), .B1 (n_207), .B2 (n_209));
INV_X1 i_1330 (.ZN (n_209), .A (n_208));
NAND2_X1 i_1329 (.ZN (n_208), .A1 (B[10]), .A2 (A[2]));
NOR2_X1 i_1328 (.ZN (n_207), .A1 (n_205), .A2 (n_206));
AOI22_X1 i_1327 (.ZN (n_206), .A1 (B[12]), .A2 (A[0]), .B1 (A[1]), .B2 (B[11]));
NOR2_X1 i_1326 (.ZN (n_205), .A1 (n_198), .A2 (n_204));
NAND2_X1 i_1325 (.ZN (n_204), .A1 (B[12]), .A2 (A[1]));
NAND2_X1 i_1324 (.ZN (n_198), .A1 (A[0]), .A2 (B[11]));
OAI21_X1 i_1323 (.ZN (n_189), .A (n_188), .B1 (n_182), .B2 (n_187));
NAND2_X1 i_1322 (.ZN (n_188), .A1 (n_182), .A2 (n_187));
OAI22_X1 i_1321 (.ZN (n_187), .A1 (n_177), .A2 (n_178), .B1 (n_175), .B2 (n_176));
NAND2_X1 i_1320 (.ZN (n_182), .A1 (n_174), .A2 (n_181));
INV_X1 i_1319 (.ZN (n_181), .A (n_167));
NAND2_X1 i_1318 (.ZN (n_178), .A1 (B[9]), .A2 (A[3]));
XNOR2_X1 i_1317 (.ZN (n_177), .A (n_175), .B (n_176));
NAND2_X1 i_1316 (.ZN (n_176), .A1 (B[8]), .A2 (A[4]));
NAND2_X1 i_1315 (.ZN (n_175), .A1 (B[7]), .A2 (A[5]));
NAND2_X1 i_1314 (.ZN (n_174), .A1 (n_168), .A2 (n_171));
NOR2_X1 i_1313 (.ZN (n_171), .A1 (n_169), .A2 (n_170));
INV_X1 i_1312 (.ZN (n_170), .A (A[6]));
INV_X1 i_1311 (.ZN (n_169), .A (B[6]));
AOI21_X1 i_1310 (.ZN (n_168), .A (n_167), .B1 (n_151), .B2 (n_166));
NOR2_X1 i_1309 (.ZN (n_167), .A1 (n_151), .A2 (n_166));
NAND2_X1 i_1308 (.ZN (n_166), .A1 (A[8]), .A2 (B[4]));
NAND2_X1 i_1307 (.ZN (n_151), .A1 (B[5]), .A2 (A[7]));
INV_X1 i_1306 (.ZN (n_150), .A (n_147));
XNOR2_X1 i_1305 (.ZN (Out[3]), .A (n_146), .B (n_149));
XNOR2_X1 i_1304 (.ZN (n_149), .A (n_148), .B (n_64));
NOR2_X1 i_1303 (.ZN (n_148), .A1 (n_66), .A2 (n_147));
NOR3_X1 i_1302 (.ZN (n_147), .A1 (n_27), .A2 (n_33), .A3 (n_29));
NAND2_X1 i_1301 (.ZN (n_146), .A1 (n_142), .A2 (n_143));
NAND2_X1 i_1300 (.ZN (n_143), .A1 (n_113), .A2 (n_140));
INV_X1 i_1299 (.ZN (n_142), .A (n_141));
NOR2_X1 i_1298 (.ZN (n_141), .A1 (n_113), .A2 (n_140));
AOI21_X1 i_1297 (.ZN (n_140), .A (n_139), .B1 (n_19), .B2 (n_21));
INV_X1 i_1296 (.ZN (n_139), .A (n_22));
XNOR2_X1 i_1295 (.ZN (n_113), .A (n_107), .B (n_25));
NOR2_X1 i_1294 (.ZN (n_107), .A1 (n_99), .A2 (n_28));
INV_X1 i_1293 (.ZN (n_99), .A (A[3]));
AOI22_X1 i_1292 (.ZN (n_66), .A1 (A[1]), .A2 (B[2]), .B1 (A[2]), .B2 (B[1]));
NAND2_X1 i_1291 (.ZN (n_64), .A1 (A[0]), .A2 (B[3]));
INV_X1 i_1290 (.ZN (n_33), .A (A[2]));
INV_X1 i_1289 (.ZN (n_31), .A (A[0]));
INV_X1 i_1288 (.ZN (n_29), .A (B[2]));
INV_X1 i_1287 (.ZN (n_28), .A (B[0]));
NAND2_X1 i_1286 (.ZN (n_27), .A1 (A[1]), .A2 (B[1]));
NAND2_X1 i_1285 (.ZN (n_26), .A1 (A[0]), .A2 (B[2]));
NOR2_X1 i_1284 (.ZN (n_25), .A1 (n_27), .A2 (n_26));
AOI21_X1 i_1283 (.ZN (n_24), .A (n_25), .B1 (n_27), .B2 (n_26));
NOR2_X1 i_1282 (.ZN (n_23), .A1 (n_33), .A2 (n_28));
NAND2_X1 i_1281 (.ZN (n_22), .A1 (n_24), .A2 (n_23));
OR2_X1 i_1280 (.ZN (n_21), .A1 (n_24), .A2 (n_23));
NAND2_X1 i_1279 (.ZN (n_20), .A1 (A[0]), .A2 (B[0]));
NOR2_X1 i_1278 (.ZN (n_19), .A1 (n_27), .A2 (n_20));
NAND2_X1 i_1277 (.ZN (n_18), .A1 (n_22), .A2 (n_21));
XNOR2_X1 i_1276 (.ZN (Out[2]), .A (n_19), .B (n_18));
AOI21_X4 i_2675 (.ZN (Out[47]), .A (n_7), .B1 (n_15), .B2 (n_17));
XNOR2_X1 i_2674 (.ZN (Out[46]), .A (n_15), .B (n_17));
XOR2_X1 i_2673 (.Z (n_17), .A (n_16), .B (n_7));
AOI21_X1 i_2672 (.ZN (n_16), .A (n_8), .B1 (n_6), .B2 (n_10));
AOI21_X1 i_2671 (.ZN (n_15), .A (n_13), .B1 (n_2597), .B2 (n_14));
AOI21_X1 i_2670 (.ZN (n_14), .A (n_1), .B1 (n_2570), .B2 (n_11));
AOI21_X1 i_1275 (.ZN (n_13), .A (n_11), .B1 (n_2580), .B2 (n_2570));
XNOR2_X1 i_2667 (.ZN (Out[45]), .A (n_5), .B (n_12));
XOR2_X1 i_2666 (.Z (n_12), .A (n_2569), .B (n_11));
XNOR2_X1 i_1274 (.ZN (n_11), .A (n_6), .B (n_10));
NOR2_X1 i_1273 (.ZN (n_10), .A1 (n_8), .A2 (n_9));
AOI22_X1 i_1272 (.ZN (n_9), .A1 (A[22]), .A2 (B[23]), .B1 (B[22]), .B2 (A[23]));
NOR2_X1 i_1271 (.ZN (n_8), .A1 (n_2517), .A2 (n_7));
NAND2_X1 i_1270 (.ZN (n_7), .A1 (B[23]), .A2 (A[23]));
OAI22_X1 i_1269 (.ZN (n_6), .A1 (n_2520), .A2 (n_2562), .B1 (n_2517), .B2 (n_2519));
AOI21_X1 i_2658 (.ZN (n_5), .A (n_1), .B1 (n_4), .B2 (n_2580));
INV_X1 i_2657 (.ZN (n_4), .A (n_2597));
XOR2_X1 i_2656 (.Z (Out[44]), .A (n_2597), .B (n_2));
NOR2_X1 i_2655 (.ZN (n_2), .A1 (n_0), .A2 (n_1));
NOR2_X1 i_2654 (.ZN (n_1), .A1 (n_2582), .A2 (n_2581));
INV_X1 i_2653 (.ZN (n_0), .A (n_2580));
AOI22_X1 i_2641 (.ZN (n_2597), .A1 (n_2578), .A2 (n_2595), .B1 (n_2594), .B2 (n_2596));
INV_X1 i_2640 (.ZN (n_2596), .A (n_2579));
XNOR2_X1 i_2639 (.ZN (Out[43]), .A (n_2578), .B (n_2595));
XNOR2_X1 i_2638 (.ZN (n_2595), .A (n_2579), .B (n_2594));
XNOR2_X1 i_2637 (.ZN (n_2594), .A (n_2592), .B (n_2583));
AOI22_X1 i_2622 (.ZN (n_2579), .A1 (n_2574), .A2 (n_2575), .B1 (n_2572), .B2 (n_2573));
OAI21_X1 i_2621 (.ZN (n_2578), .A (n_2552), .B1 (n_2577), .B2 (n_2576));
INV_X1 i_2620 (.ZN (n_2577), .A (n_2551));
XNOR2_X1 i_2619 (.ZN (Out[42]), .A (n_2553), .B (n_2576));
XNOR2_X1 i_2618 (.ZN (n_2576), .A (n_2574), .B (n_2575));
AOI21_X1 i_2617 (.ZN (n_2575), .A (n_2535), .B1 (n_2522), .B2 (n_2536));
XOR2_X1 i_2616 (.Z (n_2574), .A (n_2572), .B (n_2573));
AOI22_X1 i_2615 (.ZN (n_2573), .A1 (n_2515), .A2 (n_2357), .B1 (n_2371), .B2 (n_2360));
XNOR2_X1 i_2614 (.ZN (n_2572), .A (n_2590), .B (n_2584));
NAND2_X1 i_2595 (.ZN (n_2553), .A1 (n_2551), .A2 (n_2552));
NAND2_X1 i_2594 (.ZN (n_2552), .A1 (n_2548), .A2 (n_2550));
OR2_X1 i_2593 (.ZN (n_2551), .A1 (n_2548), .A2 (n_2550));
INV_X1 i_2592 (.ZN (n_2550), .A (n_2549));
AOI22_X1 i_2591 (.ZN (n_2549), .A1 (n_2539), .A2 (n_2542), .B1 (n_2537), .B2 (n_2538));
AOI21_X1 i_1268 (.ZN (n_2548), .A (n_2544), .B1 (n_2512), .B2 (n_2545));
XOR2_X1 i_2589 (.Z (Out[41]), .A (n_2512), .B (n_2547));
NOR2_X1 i_2588 (.ZN (n_2547), .A1 (n_2544), .A2 (n_2546));
INV_X1 i_2587 (.ZN (n_2546), .A (n_2545));
NAND2_X1 i_1267 (.ZN (n_2545), .A1 (n_2513), .A2 (n_2543));
NOR2_X1 i_1266 (.ZN (n_2544), .A1 (n_2513), .A2 (n_2543));
XOR2_X1 i_1265 (.Z (n_2543), .A (n_2539), .B (n_2542));
AOI22_X1 i_1264 (.ZN (n_2542), .A1 (n_2420), .A2 (n_2540), .B1 (n_2421), .B2 (n_2304));
INV_X1 i_1263 (.ZN (n_2540), .A (n_2406));
XOR2_X1 i_1262 (.Z (n_2539), .A (n_2537), .B (n_2538));
AOI22_X1 i_1261 (.ZN (n_2538), .A1 (n_2400), .A2 (n_2384), .B1 (n_2403), .B2 (n_2404));
XNOR2_X1 i_1260 (.ZN (n_2537), .A (n_2522), .B (n_2536));
AOI21_X1 i_1259 (.ZN (n_2536), .A (n_2535), .B1 (n_2534), .B2 (n_2527));
NOR2_X1 i_1258 (.ZN (n_2535), .A1 (n_2527), .A2 (n_2534));
OAI21_X1 i_1257 (.ZN (n_2534), .A (n_2528), .B1 (n_2526), .B2 (n_2521));
XOR2_X1 i_1256 (.Z (n_2527), .A (n_2587), .B (n_2370));
XOR2_X1 i_1255 (.Z (n_2522), .A (n_2515), .B (n_2357));
AOI21_X1 i_1254 (.ZN (n_2515), .A (n_2428), .B1 (n_2514), .B2 (n_2427));
INV_X1 i_1253 (.ZN (n_2514), .A (n_2423));
AOI22_X1 i_1252 (.ZN (n_2513), .A1 (n_2444), .A2 (n_2382), .B1 (n_2405), .B2 (n_2383));
AOI22_X1 i_1251 (.ZN (n_2512), .A1 (n_2511), .A2 (n_2510), .B1 (n_2478), .B2 (n_2509));
INV_X1 i_1250 (.ZN (n_2511), .A (n_2477));
XOR2_X1 i_2551 (.Z (Out[40]), .A (n_2477), .B (n_2510));
XOR2_X1 i_1249 (.Z (n_2510), .A (n_2478), .B (n_2509));
XNOR2_X1 i_1248 (.ZN (n_2509), .A (n_2444), .B (n_2382));
AOI22_X1 i_1247 (.ZN (n_2478), .A1 (n_2471), .A2 (n_2472), .B1 (n_2452), .B2 (n_2470));
AOI22_X1 i_1246 (.ZN (n_2477), .A1 (n_2474), .A2 (n_2475), .B1 (n_2476), .B2 (n_2473));
INV_X1 i_1245 (.ZN (n_2476), .A (n_2441));
XNOR2_X1 i_2515 (.ZN (Out[39]), .A (n_2474), .B (n_2475));
AOI22_X1 i_1244 (.ZN (n_2475), .A1 (n_2402), .A2 (n_2435), .B1 (n_2399), .B2 (n_2401));
XNOR2_X1 i_1243 (.ZN (n_2474), .A (n_2441), .B (n_2473));
XNOR2_X1 i_1242 (.ZN (n_2473), .A (n_2471), .B (n_2472));
AOI22_X1 i_1241 (.ZN (n_2472), .A1 (n_2434), .A2 (n_2416), .B1 (n_2414), .B2 (n_2415));
XOR2_X1 i_1240 (.Z (n_2471), .A (n_2452), .B (n_2470));
XOR2_X1 i_1239 (.Z (n_2470), .A (n_2417), .B (n_2407));
XNOR2_X1 i_1238 (.ZN (n_2452), .A (n_2460), .B (n_2445));
AOI21_X1 i_1237 (.ZN (n_2441), .A (n_2437), .B1 (n_2395), .B2 (n_2438));
XNOR2_X1 i_2479 (.ZN (Out[38]), .A (n_2395), .B (n_2440));
NOR2_X1 i_2478 (.ZN (n_2440), .A1 (n_2437), .A2 (n_2439));
INV_X1 i_2477 (.ZN (n_2439), .A (n_2438));
NAND2_X1 i_1236 (.ZN (n_2438), .A1 (n_2397), .A2 (n_2436));
NOR2_X1 i_1235 (.ZN (n_2437), .A1 (n_2397), .A2 (n_2436));
XOR2_X1 i_1234 (.Z (n_2436), .A (n_2402), .B (n_2435));
XNOR2_X1 i_1233 (.ZN (n_2435), .A (n_2416), .B (n_2434));
XNOR2_X1 i_1232 (.ZN (n_2434), .A (n_2462), .B (n_2461));
XOR2_X1 i_1231 (.Z (n_2416), .A (n_2414), .B (n_2415));
AOI22_X1 i_1230 (.ZN (n_2415), .A1 (n_2380), .A2 (n_2385), .B1 (n_2375), .B2 (n_2379));
XOR2_X1 i_1229 (.Z (n_2414), .A (n_2450), .B (n_2449));
XOR2_X1 i_1228 (.Z (n_2402), .A (n_2399), .B (n_2401));
AOI22_X1 i_1227 (.ZN (n_2401), .A1 (n_2359), .A2 (n_2365), .B1 (n_2303), .B2 (n_2358));
OAI22_X1 i_1226 (.ZN (n_2399), .A1 (n_2369), .A2 (n_2388), .B1 (n_2398), .B2 (n_2386));
INV_X1 i_1225 (.ZN (n_2398), .A (n_2387));
OAI22_X1 i_1224 (.ZN (n_2397), .A1 (n_2367), .A2 (n_2389), .B1 (n_2396), .B2 (n_2366));
INV_X1 i_1223 (.ZN (n_2396), .A (n_2352));
OAI22_X1 i_1222 (.ZN (n_2395), .A1 (n_2351), .A2 (n_2393), .B1 (n_2394), .B2 (n_2390));
INV_X1 i_1221 (.ZN (n_2394), .A (n_2392));
XNOR2_X1 i_2431 (.ZN (Out[37]), .A (n_2351), .B (n_2393));
XOR2_X1 i_1220 (.Z (n_2393), .A (n_2390), .B (n_2392));
AOI22_X1 i_1219 (.ZN (n_2392), .A1 (n_2299), .A2 (n_2347), .B1 (n_2391), .B2 (n_2298));
INV_X1 i_1218 (.ZN (n_2391), .A (n_2293));
XOR2_X1 i_1217 (.Z (n_2390), .A (n_2367), .B (n_2389));
XNOR2_X1 i_1216 (.ZN (n_2389), .A (n_2369), .B (n_2388));
XOR2_X1 i_1215 (.Z (n_2388), .A (n_2386), .B (n_2387));
OAI21_X1 i_1214 (.ZN (n_2387), .A (n_2344), .B1 (n_2342), .B2 (n_2334));
XNOR2_X1 i_1213 (.ZN (n_2386), .A (n_2380), .B (n_2385));
XOR2_X1 i_1212 (.Z (n_2385), .A (n_2341), .B (n_2340));
XOR2_X1 i_1211 (.Z (n_2380), .A (n_2375), .B (n_2379));
XOR2_X1 i_1210 (.Z (n_2379), .A (n_2326), .B (n_2325));
XOR2_X1 i_1209 (.Z (n_2375), .A (n_2336), .B (n_2335));
AOI22_X1 i_1208 (.ZN (n_2369), .A1 (n_2294), .A2 (n_2297), .B1 (n_2368), .B2 (n_2296));
INV_X1 i_1207 (.ZN (n_2368), .A (n_2295));
XOR2_X1 i_1206 (.Z (n_2367), .A (n_2352), .B (n_2366));
XOR2_X1 i_1205 (.Z (n_2366), .A (n_2359), .B (n_2365));
XNOR2_X1 i_1204 (.ZN (n_2365), .A (n_2467), .B (n_2466));
XNOR2_X1 i_1203 (.ZN (n_2359), .A (n_2302), .B (n_2358));
XNOR2_X1 i_1202 (.ZN (n_2358), .A (n_2455), .B (n_2454));
AOI22_X1 i_1201 (.ZN (n_2352), .A1 (n_2301), .A2 (n_2346), .B1 (n_2321), .B2 (n_2345));
AOI22_X1 i_1200 (.ZN (n_2351), .A1 (n_2290), .A2 (n_2349), .B1 (n_2350), .B2 (n_2348));
INV_X1 i_1199 (.ZN (n_2350), .A (n_2292));
XNOR2_X1 i_2386 (.ZN (Out[36]), .A (n_2290), .B (n_2349));
XNOR2_X1 i_1198 (.ZN (n_2349), .A (n_2292), .B (n_2348));
XNOR2_X1 i_1197 (.ZN (n_2348), .A (n_2299), .B (n_2347));
XNOR2_X1 i_1196 (.ZN (n_2347), .A (n_2301), .B (n_2346));
XOR2_X1 i_1195 (.Z (n_2346), .A (n_2321), .B (n_2345));
OAI21_X1 i_1194 (.ZN (n_2345), .A (n_2344), .B1 (n_2343), .B2 (n_2328));
NAND2_X1 i_1193 (.ZN (n_2344), .A1 (n_2328), .A2 (n_2343));
XOR2_X1 i_1192 (.Z (n_2343), .A (n_2334), .B (n_2342));
OAI21_X1 i_1191 (.ZN (n_2342), .A (n_2457), .B1 (n_2458), .B2 (n_2506));
XNOR2_X1 i_1190 (.ZN (n_2334), .A (n_2481), .B (n_2480));
XNOR2_X1 i_1189 (.ZN (n_2328), .A (n_2490), .B (n_2484));
XNOR2_X1 i_1188 (.ZN (n_2321), .A (n_2315), .B (n_2280));
NAND2_X1 i_1187 (.ZN (n_2315), .A1 (n_2313), .A2 (n_2281));
INV_X1 i_1186 (.ZN (n_2313), .A (n_2275));
AOI22_X1 i_1185 (.ZN (n_2301), .A1 (n_2133), .A2 (n_2075), .B1 (n_2300), .B2 (n_2134));
INV_X1 i_1184 (.ZN (n_2300), .A (n_2178));
XNOR2_X1 i_1183 (.ZN (n_2299), .A (n_2293), .B (n_2298));
XOR2_X1 i_1182 (.Z (n_2298), .A (n_2294), .B (n_2297));
XNOR2_X1 i_1181 (.ZN (n_2297), .A (n_2295), .B (n_2296));
AOI22_X1 i_1180 (.ZN (n_2296), .A1 (n_2255), .A2 (n_2262), .B1 (n_2247), .B2 (n_2254));
AOI22_X1 i_1179 (.ZN (n_2295), .A1 (n_2146), .A2 (n_2135), .B1 (n_2148), .B2 (n_2147));
AOI22_X1 i_1178 (.ZN (n_2294), .A1 (n_2238), .A2 (n_2240), .B1 (n_2232), .B2 (n_2237));
AOI22_X1 i_1177 (.ZN (n_2293), .A1 (n_2229), .A2 (n_2264), .B1 (n_2241), .B2 (n_2263));
AOI22_X1 i_1176 (.ZN (n_2292), .A1 (n_2282), .A2 (n_2291), .B1 (n_2265), .B2 (n_2074));
INV_X1 i_1175 (.ZN (n_2291), .A (n_2228));
AOI21_X1 i_1174 (.ZN (n_2290), .A (n_2289), .B1 (n_2226), .B2 (n_2286));
INV_X1 i_1173 (.ZN (n_2289), .A (n_2287));
XNOR2_X1 i_1172 (.ZN (Out[35]), .A (n_2226), .B (n_2288));
NAND2_X1 i_1171 (.ZN (n_2288), .A1 (n_2286), .A2 (n_2287));
NAND2_X1 i_1170 (.ZN (n_2287), .A1 (n_2283), .A2 (n_2285));
OR2_X1 i_1169 (.ZN (n_2286), .A1 (n_2283), .A2 (n_2285));
AOI22_X1 i_1168 (.ZN (n_2285), .A1 (n_2206), .A2 (n_2223), .B1 (n_2284), .B2 (n_2205));
INV_X1 i_1167 (.ZN (n_2284), .A (n_2171));
XOR2_X1 i_1166 (.Z (n_2283), .A (n_2228), .B (n_2282));
XOR2_X1 i_1165 (.Z (n_2282), .A (n_2265), .B (n_2074));
XNOR2_X1 i_1164 (.ZN (n_2265), .A (n_2229), .B (n_2264));
XOR2_X1 i_1163 (.Z (n_2264), .A (n_2241), .B (n_2263));
XNOR2_X1 i_1162 (.ZN (n_2263), .A (n_2255), .B (n_2262));
XNOR2_X1 i_1161 (.ZN (n_2262), .A (n_2486), .B (n_2485));
XOR2_X1 i_1160 (.Z (n_2255), .A (n_2247), .B (n_2254));
XNOR2_X1 i_1159 (.ZN (n_2254), .A (n_2501), .B (n_2500));
XNOR2_X1 i_1158 (.ZN (n_2247), .A (n_2496), .B (n_2495));
XNOR2_X1 i_1157 (.ZN (n_2241), .A (n_2238), .B (n_2240));
AOI22_X1 i_1156 (.ZN (n_2240), .A1 (n_2198), .A2 (n_2203), .B1 (n_2239), .B2 (n_2197));
INV_X1 i_1155 (.ZN (n_2239), .A (n_2193));
XOR2_X1 i_1154 (.Z (n_2238), .A (n_2232), .B (n_2237));
XNOR2_X1 i_1153 (.ZN (n_2237), .A (n_2260), .B (n_2261));
AOI22_X1 i_1152 (.ZN (n_2232), .A1 (n_2230), .A2 (n_2195), .B1 (n_2210), .B2 (n_2231));
INV_X1 i_1151 (.ZN (n_2231), .A (n_2196));
INV_X1 i_1150 (.ZN (n_2230), .A (n_2216));
AOI22_X1 i_1149 (.ZN (n_2229), .A1 (n_2191), .A2 (n_2204), .B1 (n_2190), .B2 (n_2189));
AOI22_X1 i_1148 (.ZN (n_2228), .A1 (n_2227), .A2 (n_2222), .B1 (n_2221), .B2 (n_2219));
INV_X1 i_1147 (.ZN (n_2227), .A (n_2208));
AOI22_X1 i_1146 (.ZN (n_2226), .A1 (n_2169), .A2 (n_2225), .B1 (n_2224), .B2 (n_2170));
XNOR2_X1 i_1145 (.ZN (Out[34]), .A (n_2169), .B (n_2225));
XOR2_X1 i_1144 (.Z (n_2225), .A (n_2170), .B (n_2224));
XOR2_X1 i_1143 (.Z (n_2224), .A (n_2206), .B (n_2223));
XNOR2_X1 i_1142 (.ZN (n_2223), .A (n_2208), .B (n_2222));
XOR2_X1 i_1141 (.Z (n_2222), .A (n_2219), .B (n_2221));
AOI22_X1 i_1140 (.ZN (n_2221), .A1 (n_2157), .A2 (n_2220), .B1 (n_2155), .B2 (n_2156));
INV_X1 i_1139 (.ZN (n_2220), .A (n_2159));
XOR2_X1 i_1138 (.Z (n_2219), .A (n_2085), .B (n_2076));
AOI22_X1 i_1137 (.ZN (n_2208), .A1 (n_2139), .A2 (n_2207), .B1 (n_2121), .B2 (n_2138));
INV_X1 i_1136 (.ZN (n_2207), .A (n_2103));
XNOR2_X1 i_1135 (.ZN (n_2206), .A (n_2171), .B (n_2205));
XOR2_X1 i_1134 (.Z (n_2205), .A (n_2191), .B (n_2204));
XNOR2_X1 i_1133 (.ZN (n_2204), .A (n_2198), .B (n_2203));
XOR2_X1 i_1132 (.Z (n_2203), .A (n_2253), .B (n_2256));
XNOR2_X1 i_1131 (.ZN (n_2198), .A (n_2193), .B (n_2197));
XOR2_X1 i_1130 (.Z (n_2197), .A (n_2246), .B (n_2248));
AOI22_X1 i_1129 (.ZN (n_2193), .A1 (n_2107), .A2 (n_2087), .B1 (n_2192), .B2 (n_2109));
INV_X1 i_1128 (.ZN (n_2192), .A (n_2110));
XOR2_X1 i_1127 (.Z (n_2191), .A (n_2189), .B (n_2190));
AOI22_X1 i_1126 (.ZN (n_2190), .A1 (n_2113), .A2 (n_2120), .B1 (n_2106), .B2 (n_2112));
XNOR2_X1 i_1125 (.ZN (n_2189), .A (n_2194), .B (n_2179));
AOI22_X1 i_1124 (.ZN (n_2171), .A1 (n_2073), .A2 (n_2161), .B1 (n_2144), .B2 (n_2160));
AOI22_X1 i_1123 (.ZN (n_2170), .A1 (n_2141), .A2 (n_2162), .B1 (n_2140), .B2 (n_2101));
AOI21_X1 i_1122 (.ZN (n_2169), .A (n_2168), .B1 (n_2099), .B2 (n_2165));
INV_X1 i_1121 (.ZN (n_2168), .A (n_2166));
XNOR2_X1 i_1120 (.ZN (Out[33]), .A (n_2099), .B (n_2167));
NAND2_X1 i_1119 (.ZN (n_2167), .A1 (n_2165), .A2 (n_2166));
NAND2_X1 i_1118 (.ZN (n_2166), .A1 (n_2163), .A2 (n_2164));
OR2_X1 i_1117 (.ZN (n_2165), .A1 (n_2163), .A2 (n_2164));
AOI22_X1 i_1116 (.ZN (n_2164), .A1 (n_2093), .A2 (n_2090), .B1 (n_2089), .B2 (n_2051));
XOR2_X1 i_1115 (.Z (n_2163), .A (n_2141), .B (n_2162));
XNOR2_X1 i_1114 (.ZN (n_2162), .A (n_2073), .B (n_2161));
XOR2_X1 i_1113 (.Z (n_2161), .A (n_2144), .B (n_2160));
XOR2_X1 i_1112 (.Z (n_2160), .A (n_2157), .B (n_2159));
AOI22_X1 i_1111 (.ZN (n_2159), .A1 (n_1991), .A2 (n_2038), .B1 (n_2158), .B2 (n_1990));
INV_X1 i_1110 (.ZN (n_2158), .A (n_1984));
XOR2_X1 i_1109 (.Z (n_2157), .A (n_2155), .B (n_2156));
AOI22_X1 i_1108 (.ZN (n_2156), .A1 (n_1976), .A2 (n_1981), .B1 (n_1962), .B2 (n_1975));
XOR2_X1 i_1107 (.Z (n_2155), .A (n_2086), .B (n_2111));
AOI22_X1 i_1106 (.ZN (n_2144), .A1 (n_2028), .A2 (n_2029), .B1 (n_2027), .B2 (n_1894));
XOR2_X1 i_1105 (.Z (n_2141), .A (n_2101), .B (n_2140));
XOR2_X1 i_1104 (.Z (n_2140), .A (n_2103), .B (n_2139));
XOR2_X1 i_1103 (.Z (n_2139), .A (n_2121), .B (n_2138));
XOR2_X1 i_1102 (.Z (n_2138), .A (n_2081), .B (n_2080));
XNOR2_X1 i_1101 (.ZN (n_2121), .A (n_2113), .B (n_2120));
XOR2_X1 i_1100 (.Z (n_2120), .A (n_2217), .B (n_2218));
XOR2_X1 i_1099 (.Z (n_2113), .A (n_2106), .B (n_2112));
XOR2_X1 i_1098 (.Z (n_2112), .A (n_2212), .B (n_2211));
OAI22_X1 i_1097 (.ZN (n_2106), .A1 (n_2032), .A2 (n_2035), .B1 (n_2104), .B2 (n_2105));
INV_X1 i_1096 (.ZN (n_2105), .A (n_2034));
INV_X1 i_1095 (.ZN (n_2104), .A (n_2033));
AOI22_X1 i_1094 (.ZN (n_2103), .A1 (n_2043), .A2 (n_2102), .B1 (n_2036), .B2 (n_2042));
INV_X1 i_1093 (.ZN (n_2102), .A (n_2044));
AOI21_X1 i_1092 (.ZN (n_2101), .A (n_2100), .B1 (n_2030), .B2 (n_2048));
INV_X1 i_1091 (.ZN (n_2100), .A (n_2049));
AOI21_X1 i_1090 (.ZN (n_2099), .A (n_2095), .B1 (n_2023), .B2 (n_2096));
XNOR2_X1 i_1089 (.ZN (Out[32]), .A (n_2023), .B (n_2098));
NOR2_X1 i_1088 (.ZN (n_2098), .A1 (n_2095), .A2 (n_2097));
INV_X1 i_1087 (.ZN (n_2097), .A (n_2096));
NAND2_X1 i_1086 (.ZN (n_2096), .A1 (n_2024), .A2 (n_2094));
NOR2_X1 i_1085 (.ZN (n_2095), .A1 (n_2024), .A2 (n_2094));
XNOR2_X1 i_1084 (.ZN (n_2094), .A (n_2090), .B (n_2093));
AOI22_X1 i_1083 (.ZN (n_2093), .A1 (n_1971), .A2 (n_2091), .B1 (n_1968), .B2 (n_2092));
INV_X1 i_1082 (.ZN (n_2092), .A (n_1970));
INV_X1 i_1081 (.ZN (n_2091), .A (n_1972));
XOR2_X1 i_1080 (.Z (n_2090), .A (n_2051), .B (n_2089));
XOR2_X1 i_1079 (.Z (n_2089), .A (n_2068), .B (n_2071));
XNOR2_X1 i_1078 (.ZN (n_2051), .A (n_2030), .B (n_2050));
NAND2_X1 i_1077 (.ZN (n_2050), .A1 (n_2048), .A2 (n_2049));
NAND2_X1 i_1076 (.ZN (n_2049), .A1 (n_2045), .A2 (n_2047));
OR2_X1 i_1075 (.ZN (n_2048), .A1 (n_2045), .A2 (n_2047));
OAI21_X1 i_1074 (.ZN (n_2047), .A (n_2001), .B1 (n_2015), .B2 (n_2046));
INV_X1 i_1073 (.ZN (n_2046), .A (n_2000));
XNOR2_X1 i_1072 (.ZN (n_2045), .A (n_2043), .B (n_2044));
AOI22_X1 i_1071 (.ZN (n_2044), .A1 (n_1994), .A2 (n_1998), .B1 (n_1989), .B2 (n_1993));
XOR2_X1 i_1070 (.Z (n_2043), .A (n_2036), .B (n_2042));
XNOR2_X1 i_1069 (.ZN (n_2042), .A (n_2125), .B (n_2118));
XNOR2_X1 i_1068 (.ZN (n_2036), .A (n_2032), .B (n_2035));
XNOR2_X1 i_1067 (.ZN (n_2035), .A (n_2033), .B (n_2034));
OAI22_X1 i_1066 (.ZN (n_2034), .A1 (n_2004), .A2 (n_2005), .B1 (n_1840), .B2 (n_2132));
OAI22_X1 i_1065 (.ZN (n_2033), .A1 (n_1996), .A2 (n_1997), .B1 (n_1929), .B2 (n_1995));
AOI22_X1 i_1064 (.ZN (n_2032), .A1 (n_2012), .A2 (n_2013), .B1 (n_2010), .B2 (n_2031));
INV_X1 i_1063 (.ZN (n_2031), .A (n_2011));
XNOR2_X1 i_1062 (.ZN (n_2030), .A (n_2028), .B (n_2029));
AOI22_X1 i_1061 (.ZN (n_2029), .A1 (n_2014), .A2 (n_2009), .B1 (n_2008), .B2 (n_2006));
XOR2_X1 i_1060 (.Z (n_2028), .A (n_1894), .B (n_2027));
OAI21_X1 i_1059 (.ZN (n_2027), .A (n_2060), .B1 (n_2053), .B2 (n_2052));
AOI22_X1 i_1058 (.ZN (n_2024), .A1 (n_2017), .A2 (n_2018), .B1 (n_1973), .B2 (n_2016));
OAI21_X1 i_1057 (.ZN (n_2023), .A (n_2022), .B1 (n_2020), .B2 (n_2019));
OAI21_X1 i_1056 (.ZN (Out[31]), .A (n_2022), .B1 (n_1950), .B2 (n_2021));
NAND2_X1 i_1055 (.ZN (n_2022), .A1 (n_1950), .A2 (n_2021));
XOR2_X1 i_1054 (.Z (n_2021), .A (n_2019), .B (n_2020));
AOI22_X1 i_1053 (.ZN (n_2020), .A1 (n_1901), .A2 (n_1944), .B1 (n_1867), .B2 (n_1900));
XNOR2_X1 i_1052 (.ZN (n_2019), .A (n_2017), .B (n_2018));
OAI22_X1 i_1051 (.ZN (n_2018), .A1 (n_1902), .A2 (n_1943), .B1 (n_1904), .B2 (n_1942));
XOR2_X1 i_1050 (.Z (n_2017), .A (n_1973), .B (n_2016));
XOR2_X1 i_1049 (.Z (n_2016), .A (n_2002), .B (n_2015));
XNOR2_X1 i_1048 (.ZN (n_2015), .A (n_2009), .B (n_2014));
XNOR2_X1 i_1047 (.ZN (n_2014), .A (n_2012), .B (n_2013));
AOI21_X1 i_1046 (.ZN (n_2013), .A (n_1837), .B1 (n_1838), .B2 (n_1841));
XNOR2_X1 i_1045 (.ZN (n_2012), .A (n_2010), .B (n_2011));
AOI21_X1 i_1044 (.ZN (n_2011), .A (n_1928), .B1 (n_1926), .B2 (n_1925));
OAI33_X1 i_1043 (.ZN (n_2010), .A1 (n_1912), .A2 (n_558), .A3 (n_560), .B1 (n_1848)
    , .B2 (n_256), .B3 (n_1232));
XOR2_X1 i_1042 (.Z (n_2009), .A (n_2006), .B (n_2008));
AOI22_X1 i_1041 (.ZN (n_2008), .A1 (n_1823), .A2 (n_1814), .B1 (n_2007), .B2 (n_1815));
INV_X1 i_1040 (.ZN (n_2007), .A (n_1821));
XNOR2_X1 i_1039 (.ZN (n_2006), .A (n_2004), .B (n_2005));
NAND2_X1 i_1038 (.ZN (n_2005), .A1 (A[8]), .A2 (B[23]));
XNOR2_X1 i_1037 (.ZN (n_2004), .A (n_1840), .B (n_2132));
NAND2_X1 i_1036 (.ZN (n_2002), .A1 (n_2000), .A2 (n_2001));
NAND2_X1 i_1035 (.ZN (n_2001), .A1 (n_1983), .A2 (n_1999));
OR2_X1 i_1034 (.ZN (n_2000), .A1 (n_1983), .A2 (n_1999));
XOR2_X1 i_1033 (.Z (n_1999), .A (n_1994), .B (n_1998));
XNOR2_X1 i_1032 (.ZN (n_1998), .A (n_1996), .B (n_1997));
NAND2_X1 i_1031 (.ZN (n_1997), .A1 (A[11]), .A2 (B[20]));
XNOR2_X1 i_1030 (.ZN (n_1996), .A (n_1929), .B (n_1995));
NAND2_X1 i_1029 (.ZN (n_1995), .A1 (A[13]), .A2 (B[18]));
XOR2_X1 i_1028 (.Z (n_1994), .A (n_1989), .B (n_1993));
XNOR2_X1 i_1027 (.ZN (n_1993), .A (n_2131), .B (n_2130));
XNOR2_X1 i_1026 (.ZN (n_1989), .A (n_2119), .B (n_1964));
XOR2_X1 i_1025 (.Z (n_1983), .A (n_1895), .B (n_1930));
XOR2_X1 i_1024 (.Z (n_1973), .A (n_1971), .B (n_1972));
AOI22_X1 i_1023 (.ZN (n_1972), .A1 (n_1793), .A2 (n_1899), .B1 (n_1812), .B2 (n_1794));
XNOR2_X1 i_1022 (.ZN (n_1971), .A (n_1968), .B (n_1970));
AOI21_X1 i_1021 (.ZN (n_1970), .A (n_1969), .B1 (n_1892), .B2 (n_1939));
INV_X1 i_1020 (.ZN (n_1969), .A (n_1938));
XOR2_X1 i_1019 (.Z (n_1968), .A (n_2064), .B (n_2066));
OAI21_X1 i_1018 (.ZN (n_1950), .A (n_1947), .B1 (n_1863), .B2 (n_1949));
INV_X1 i_1017 (.ZN (n_1949), .A (n_1946));
XNOR2_X1 i_1016 (.ZN (Out[30]), .A (n_1863), .B (n_1948));
NAND2_X1 i_1015 (.ZN (n_1948), .A1 (n_1946), .A2 (n_1947));
OR2_X1 i_1014 (.ZN (n_1947), .A1 (n_1945), .A2 (n_1866));
NAND2_X1 i_1013 (.ZN (n_1946), .A1 (n_1866), .A2 (n_1945));
XNOR2_X1 i_1012 (.ZN (n_1945), .A (n_1901), .B (n_1944));
XOR2_X1 i_1011 (.Z (n_1944), .A (n_1902), .B (n_1943));
XNOR2_X1 i_1010 (.ZN (n_1943), .A (n_1904), .B (n_1942));
XNOR2_X1 i_1009 (.ZN (n_1942), .A (n_1940), .B (n_1892));
NAND2_X1 i_1008 (.ZN (n_1940), .A1 (n_1938), .A2 (n_1939));
NAND2_X1 i_1007 (.ZN (n_1939), .A1 (n_1919), .A2 (n_1937));
OR2_X1 i_1006 (.ZN (n_1938), .A1 (n_1919), .A2 (n_1937));
XOR2_X1 i_1005 (.Z (n_1937), .A (n_1914), .B (n_1910));
XNOR2_X1 i_1004 (.ZN (n_1919), .A (n_1935), .B (n_1931));
AOI22_X1 i_1003 (.ZN (n_1904), .A1 (n_1836), .A2 (n_1854), .B1 (n_1535), .B2 (n_1903));
INV_X1 i_1002 (.ZN (n_1903), .A (n_1835));
AOI22_X1 i_1001 (.ZN (n_1902), .A1 (n_1799), .A2 (n_1817), .B1 (n_1718), .B2 (n_1798));
XOR2_X1 i_1000 (.Z (n_1901), .A (n_1867), .B (n_1900));
XNOR2_X1 i_999 (.ZN (n_1900), .A (n_1793), .B (n_1899));
AOI22_X1 i_998 (.ZN (n_1899), .A1 (n_1898), .A2 (n_1816), .B1 (n_1719), .B2 (n_1804));
INV_X1 i_997 (.ZN (n_1898), .A (n_1802));
AOI22_X1 i_996 (.ZN (n_1867), .A1 (n_1856), .A2 (n_1857), .B1 (n_1820), .B2 (n_1855));
INV_X1 i_995 (.ZN (n_1866), .A (n_1865));
AOI22_X1 i_994 (.ZN (n_1865), .A1 (n_1819), .A2 (n_1858), .B1 (n_1864), .B2 (n_1818));
INV_X1 i_993 (.ZN (n_1864), .A (n_1781));
AOI22_X1 i_992 (.ZN (n_1863), .A1 (n_1780), .A2 (n_1862), .B1 (n_1859), .B2 (n_1861));
XNOR2_X1 i_991 (.ZN (Out[29]), .A (n_1780), .B (n_1862));
XOR2_X1 i_990 (.Z (n_1862), .A (n_1859), .B (n_1861));
AOI22_X1 i_989 (.ZN (n_1861), .A1 (n_1751), .A2 (n_1778), .B1 (n_1860), .B2 (n_1750));
INV_X1 i_988 (.ZN (n_1860), .A (n_1697));
XNOR2_X1 i_987 (.ZN (n_1859), .A (n_1819), .B (n_1858));
XOR2_X1 i_986 (.Z (n_1858), .A (n_1856), .B (n_1857));
AOI22_X1 i_985 (.ZN (n_1857), .A1 (n_1727), .A2 (n_1749), .B1 (n_1729), .B2 (n_1748));
XOR2_X1 i_984 (.Z (n_1856), .A (n_1820), .B (n_1855));
XNOR2_X1 i_983 (.ZN (n_1855), .A (n_1836), .B (n_1854));
XOR2_X1 i_982 (.Z (n_1854), .A (n_1806), .B (n_1805));
XNOR2_X1 i_981 (.ZN (n_1836), .A (n_1535), .B (n_1835));
AOI22_X1 i_980 (.ZN (n_1835), .A1 (n_1742), .A2 (n_1747), .B1 (n_1735), .B2 (n_1741));
AOI22_X1 i_979 (.ZN (n_1820), .A1 (n_1766), .A2 (n_1772), .B1 (n_1752), .B2 (n_1765));
XNOR2_X1 i_978 (.ZN (n_1819), .A (n_1781), .B (n_1818));
XNOR2_X1 i_977 (.ZN (n_1818), .A (n_1799), .B (n_1817));
XNOR2_X1 i_976 (.ZN (n_1817), .A (n_1802), .B (n_1816));
XOR2_X1 i_975 (.Z (n_1816), .A (n_1804), .B (n_1719));
AOI22_X1 i_974 (.ZN (n_1804), .A1 (n_1759), .A2 (n_1764), .B1 (n_1803), .B2 (n_1758));
INV_X1 i_973 (.ZN (n_1803), .A (n_1753));
AOI22_X1 i_972 (.ZN (n_1802), .A1 (n_1800), .A2 (n_1771), .B1 (n_1801), .B2 (n_1770));
INV_X1 i_971 (.ZN (n_1801), .A (n_1769));
INV_X1 i_970 (.ZN (n_1800), .A (n_1768));
XOR2_X1 i_969 (.Z (n_1799), .A (n_1718), .B (n_1798));
OAI21_X1 i_968 (.ZN (n_1798), .A (n_1891), .B1 (n_1889), .B2 (n_1890));
AOI22_X1 i_967 (.ZN (n_1781), .A1 (n_1775), .A2 (n_1777), .B1 (n_1773), .B2 (n_1774));
OAI22_X1 i_966 (.ZN (n_1780), .A1 (n_1696), .A2 (n_1779), .B1 (n_1694), .B2 (n_1695));
XNOR2_X1 i_965 (.ZN (Out[28]), .A (n_1696), .B (n_1779));
XOR2_X1 i_964 (.Z (n_1779), .A (n_1751), .B (n_1778));
XOR2_X1 i_963 (.Z (n_1778), .A (n_1775), .B (n_1777));
AOI22_X1 i_962 (.ZN (n_1777), .A1 (n_1642), .A2 (n_1776), .B1 (n_1618), .B2 (n_1641));
INV_X1 i_961 (.ZN (n_1776), .A (n_1644));
XOR2_X1 i_960 (.Z (n_1775), .A (n_1773), .B (n_1774));
AOI22_X1 i_959 (.ZN (n_1774), .A1 (n_1667), .A2 (n_1683), .B1 (n_1444), .B2 (n_1666));
XNOR2_X1 i_958 (.ZN (n_1773), .A (n_1766), .B (n_1772));
XNOR2_X1 i_957 (.ZN (n_1772), .A (n_1768), .B (n_1771));
XNOR2_X1 i_956 (.ZN (n_1771), .A (n_1769), .B (n_1770));
OAI21_X1 i_955 (.ZN (n_1770), .A (n_1664), .B1 (n_1656), .B2 (n_1651));
AOI22_X1 i_954 (.ZN (n_1769), .A1 (n_1633), .A2 (n_1637), .B1 (n_1625), .B2 (n_1632));
AOI22_X1 i_953 (.ZN (n_1768), .A1 (n_1672), .A2 (n_1678), .B1 (n_1668), .B2 (n_1767));
INV_X1 i_952 (.ZN (n_1767), .A (n_1671));
XOR2_X1 i_951 (.Z (n_1766), .A (n_1752), .B (n_1765));
XNOR2_X1 i_950 (.ZN (n_1765), .A (n_1759), .B (n_1764));
XOR2_X1 i_949 (.Z (n_1764), .A (n_1877), .B (n_1878));
XNOR2_X1 i_948 (.ZN (n_1759), .A (n_1753), .B (n_1758));
XNOR2_X1 i_947 (.ZN (n_1758), .A (n_1756), .B (n_1882));
NAND2_X1 i_946 (.ZN (n_1756), .A1 (n_1893), .A2 (n_1880));
AOI22_X1 i_945 (.ZN (n_1753), .A1 (n_1675), .A2 (n_1677), .B1 (n_1673), .B2 (n_1674));
AOI22_X1 i_944 (.ZN (n_1752), .A1 (n_1679), .A2 (n_1682), .B1 (n_1681), .B2 (n_1680));
XNOR2_X1 i_943 (.ZN (n_1751), .A (n_1697), .B (n_1750));
XNOR2_X1 i_942 (.ZN (n_1750), .A (n_1727), .B (n_1749));
XOR2_X1 i_941 (.Z (n_1749), .A (n_1729), .B (n_1748));
XOR2_X1 i_940 (.Z (n_1748), .A (n_1742), .B (n_1747));
XOR2_X1 i_939 (.Z (n_1747), .A (n_1784), .B (n_1760));
XOR2_X1 i_938 (.Z (n_1742), .A (n_1735), .B (n_1741));
XNOR2_X1 i_937 (.ZN (n_1741), .A (n_1825), .B (n_1573));
XNOR2_X1 i_936 (.ZN (n_1735), .A (n_1734), .B (n_1730));
AOI22_X1 i_935 (.ZN (n_1729), .A1 (n_1448), .A2 (n_1639), .B1 (n_1619), .B2 (n_1638));
XNOR2_X1 i_934 (.ZN (n_1727), .A (n_1662), .B (n_1717));
AOI22_X1 i_933 (.ZN (n_1697), .A1 (n_1687), .A2 (n_1689), .B1 (n_1684), .B2 (n_1686));
XNOR2_X1 i_932 (.ZN (n_1696), .A (n_1694), .B (n_1695));
OAI22_X1 i_931 (.ZN (n_1695), .A1 (n_1646), .A2 (n_1690), .B1 (n_1600), .B2 (n_1645));
AOI22_X1 i_930 (.ZN (n_1694), .A1 (n_1598), .A2 (n_1693), .B1 (n_1691), .B2 (n_1692));
XNOR2_X1 i_929 (.ZN (Out[27]), .A (n_1598), .B (n_1693));
XOR2_X1 i_928 (.Z (n_1693), .A (n_1691), .B (n_1692));
AOI22_X1 i_927 (.ZN (n_1692), .A1 (n_1517), .A2 (n_1595), .B1 (n_1516), .B2 (n_1514));
XNOR2_X1 i_926 (.ZN (n_1691), .A (n_1646), .B (n_1690));
XNOR2_X1 i_925 (.ZN (n_1690), .A (n_1687), .B (n_1689));
AOI22_X1 i_924 (.ZN (n_1689), .A1 (n_1512), .A2 (n_1688), .B1 (n_1510), .B2 (n_1511));
INV_X1 i_923 (.ZN (n_1688), .A (n_1513));
XOR2_X1 i_922 (.Z (n_1687), .A (n_1684), .B (n_1686));
AOI22_X1 i_921 (.ZN (n_1686), .A1 (n_1547), .A2 (n_1685), .B1 (n_1536), .B2 (n_1546));
INV_X1 i_920 (.ZN (n_1685), .A (n_1549));
XNOR2_X1 i_919 (.ZN (n_1684), .A (n_1667), .B (n_1683));
XNOR2_X1 i_918 (.ZN (n_1683), .A (n_1679), .B (n_1682));
XOR2_X1 i_917 (.Z (n_1682), .A (n_1680), .B (n_1681));
AOI22_X1 i_916 (.ZN (n_1681), .A1 (n_1585), .A2 (n_1591), .B1 (n_1584), .B2 (n_1578));
AOI22_X1 i_915 (.ZN (n_1680), .A1 (n_1565), .A2 (n_1570), .B1 (n_1556), .B2 (n_1564));
XNOR2_X1 i_914 (.ZN (n_1679), .A (n_1672), .B (n_1678));
XNOR2_X1 i_913 (.ZN (n_1678), .A (n_1675), .B (n_1677));
NOR2_X1 i_912 (.ZN (n_1677), .A1 (n_1029), .A2 (n_1881));
XOR2_X1 i_911 (.Z (n_1675), .A (n_1673), .B (n_1674));
NOR2_X1 i_910 (.ZN (n_1674), .A1 (n_340), .A2 (n_1792));
OAI21_X1 i_909 (.ZN (n_1673), .A (n_1581), .B1 (n_1583), .B2 (n_1318));
XNOR2_X1 i_908 (.ZN (n_1672), .A (n_1668), .B (n_1671));
OAI22_X1 i_907 (.ZN (n_1671), .A1 (n_1540), .A2 (n_1669), .B1 (n_1670), .B2 (n_1539));
INV_X1 i_906 (.ZN (n_1670), .A (n_1538));
INV_X1 i_905 (.ZN (n_1669), .A (n_1541));
AOI22_X1 i_904 (.ZN (n_1668), .A1 (n_1509), .A2 (n_1503), .B1 (n_1521), .B2 (n_1525));
XOR2_X1 i_903 (.Z (n_1667), .A (n_1444), .B (n_1666));
AOI21_X1 i_902 (.ZN (n_1666), .A (n_1665), .B1 (n_1663), .B2 (n_1657));
INV_X1 i_901 (.ZN (n_1665), .A (n_1664));
OR2_X1 i_900 (.ZN (n_1664), .A1 (n_1657), .A2 (n_1663));
XOR2_X1 i_899 (.Z (n_1663), .A (n_1739), .B (n_1738));
XNOR2_X1 i_898 (.ZN (n_1657), .A (n_1651), .B (n_1656));
XNOR2_X1 i_897 (.ZN (n_1656), .A (n_1762), .B (n_1648));
XOR2_X1 i_896 (.Z (n_1651), .A (n_1788), .B (n_1787));
XNOR2_X1 i_895 (.ZN (n_1646), .A (n_1600), .B (n_1645));
XNOR2_X1 i_894 (.ZN (n_1645), .A (n_1642), .B (n_1644));
AOI22_X1 i_893 (.ZN (n_1644), .A1 (n_1572), .A2 (n_1592), .B1 (n_1643), .B2 (n_1571));
INV_X1 i_892 (.ZN (n_1643), .A (n_1552));
XOR2_X1 i_891 (.Z (n_1642), .A (n_1618), .B (n_1641));
XOR2_X1 i_890 (.Z (n_1641), .A (n_1639), .B (n_1449));
XOR2_X1 i_889 (.Z (n_1639), .A (n_1619), .B (n_1638));
XNOR2_X1 i_888 (.ZN (n_1638), .A (n_1633), .B (n_1637));
XNOR2_X1 i_887 (.ZN (n_1637), .A (n_1612), .B (n_1611));
XOR2_X1 i_886 (.Z (n_1633), .A (n_1625), .B (n_1632));
OAI21_X1 i_885 (.ZN (n_1632), .A (n_1745), .B1 (n_1746), .B2 (n_1791));
XNOR2_X1 i_884 (.ZN (n_1625), .A (n_1731), .B (n_1710));
OAI21_X1 i_883 (.ZN (n_1619), .A (n_1543), .B1 (n_1544), .B2 (n_1545));
XNOR2_X1 i_882 (.ZN (n_1618), .A (n_1655), .B (n_1658));
AOI22_X1 i_881 (.ZN (n_1600), .A1 (n_1599), .A2 (n_1594), .B1 (n_1550), .B2 (n_1593));
INV_X1 i_880 (.ZN (n_1599), .A (n_1520));
OAI22_X1 i_879 (.ZN (n_1598), .A1 (n_1498), .A2 (n_1597), .B1 (n_1500), .B2 (n_1596));
XNOR2_X1 i_878 (.ZN (Out[26]), .A (n_1498), .B (n_1597));
XNOR2_X1 i_877 (.ZN (n_1597), .A (n_1500), .B (n_1596));
XOR2_X1 i_876 (.Z (n_1596), .A (n_1517), .B (n_1595));
XNOR2_X1 i_875 (.ZN (n_1595), .A (n_1520), .B (n_1594));
XOR2_X1 i_874 (.Z (n_1594), .A (n_1550), .B (n_1593));
XNOR2_X1 i_873 (.ZN (n_1593), .A (n_1572), .B (n_1592));
XOR2_X1 i_872 (.Z (n_1592), .A (n_1585), .B (n_1591));
XNOR2_X1 i_871 (.ZN (n_1591), .A (n_1627), .B (n_1626));
XOR2_X1 i_870 (.Z (n_1585), .A (n_1578), .B (n_1584));
XNOR2_X1 i_869 (.ZN (n_1584), .A (n_1583), .B (n_1318));
NAND2_X1 i_868 (.ZN (n_1583), .A1 (n_1581), .A2 (n_1582));
OAI22_X1 i_867 (.ZN (n_1582), .A1 (n_1029), .A2 (n_1317), .B1 (n_424), .B2 (n_1792));
NAND3_X1 i_866 (.ZN (n_1581), .A1 (n_1786), .A2 (B[3]), .A3 (A[21]));
XOR2_X1 i_865 (.Z (n_1578), .A (n_1636), .B (n_1635));
XNOR2_X1 i_864 (.ZN (n_1572), .A (n_1552), .B (n_1571));
XOR2_X1 i_863 (.Z (n_1571), .A (n_1565), .B (n_1570));
XOR2_X1 i_862 (.Z (n_1570), .A (n_1587), .B (n_1508));
XOR2_X1 i_861 (.Z (n_1565), .A (n_1556), .B (n_1564));
OAI21_X1 i_860 (.ZN (n_1564), .A (n_1601), .B1 (n_1604), .B2 (n_1602));
XNOR2_X1 i_859 (.ZN (n_1556), .A (n_1616), .B (n_1615));
AOI22_X1 i_858 (.ZN (n_1552), .A1 (n_1408), .A2 (n_1416), .B1 (n_1551), .B2 (n_1407));
INV_X1 i_857 (.ZN (n_1551), .A (n_1401));
XOR2_X1 i_856 (.Z (n_1550), .A (n_1547), .B (n_1549));
AOI22_X1 i_855 (.ZN (n_1549), .A1 (n_1487), .A2 (n_1488), .B1 (n_1548), .B2 (n_1486));
INV_X1 i_854 (.ZN (n_1548), .A (n_1475));
XOR2_X1 i_853 (.Z (n_1547), .A (n_1536), .B (n_1546));
XNOR2_X1 i_852 (.ZN (n_1546), .A (n_1544), .B (n_1545));
OAI22_X1 i_851 (.ZN (n_1545), .A1 (n_1440), .A2 (n_1445), .B1 (n_1435), .B2 (n_1439));
OAI21_X1 i_850 (.ZN (n_1544), .A (n_1543), .B1 (n_1537), .B2 (n_1542));
NAND2_X1 i_849 (.ZN (n_1543), .A1 (n_1537), .A2 (n_1542));
XNOR2_X1 i_848 (.ZN (n_1542), .A (n_1540), .B (n_1541));
OAI22_X1 i_847 (.ZN (n_1541), .A1 (n_1437), .A2 (n_1438), .B1 (n_1344), .B2 (n_1631));
XOR2_X1 i_846 (.Z (n_1540), .A (n_1538), .B (n_1539));
AOI21_X1 i_845 (.ZN (n_1539), .A (n_1319), .B1 (n_1321), .B2 (n_1323));
OAI22_X1 i_844 (.ZN (n_1538), .A1 (n_1433), .A2 (n_1434), .B1 (n_1375), .B2 (n_1432));
AOI22_X1 i_843 (.ZN (n_1537), .A1 (n_1458), .A2 (n_1463), .B1 (n_1451), .B2 (n_1457));
XNOR2_X1 i_842 (.ZN (n_1536), .A (n_1502), .B (n_1450));
AOI22_X1 i_841 (.ZN (n_1520), .A1 (n_1518), .A2 (n_1490), .B1 (n_1519), .B2 (n_1489));
INV_X1 i_840 (.ZN (n_1519), .A (n_1473));
INV_X1 i_839 (.ZN (n_1518), .A (n_1492));
XOR2_X1 i_838 (.Z (n_1517), .A (n_1514), .B (n_1516));
OAI22_X1 i_837 (.ZN (n_1516), .A1 (n_1468), .A2 (n_1470), .B1 (n_1430), .B2 (n_1515));
INV_X1 i_836 (.ZN (n_1515), .A (n_1467));
XOR2_X1 i_835 (.Z (n_1514), .A (n_1512), .B (n_1513));
AOI22_X1 i_834 (.ZN (n_1513), .A1 (n_1428), .A2 (n_1429), .B1 (n_1417), .B2 (n_1427));
XOR2_X1 i_833 (.Z (n_1512), .A (n_1510), .B (n_1511));
OAI21_X1 i_832 (.ZN (n_1511), .A (n_1466), .B1 (n_1446), .B2 (n_1464));
XNOR2_X1 i_831 (.ZN (n_1510), .A (n_1413), .B (n_1443));
AOI22_X1 i_830 (.ZN (n_1500), .A1 (n_1494), .A2 (n_1499), .B1 (n_1471), .B2 (n_1493));
INV_X1 i_829 (.ZN (n_1499), .A (n_1495));
AOI21_X1 i_828 (.ZN (n_1498), .A (n_1496), .B1 (n_1399), .B2 (n_1497));
XNOR2_X1 i_827 (.ZN (Out[25]), .A (n_1399), .B (n_1497));
XNOR2_X1 i_826 (.ZN (n_1497), .A (n_1496), .B (n_1397));
XNOR2_X1 i_825 (.ZN (n_1496), .A (n_1494), .B (n_1495));
AOI22_X1 i_824 (.ZN (n_1495), .A1 (n_1313), .A2 (n_1393), .B1 (n_1312), .B2 (n_1310));
XOR2_X1 i_823 (.Z (n_1494), .A (n_1471), .B (n_1493));
XOR2_X1 i_822 (.Z (n_1493), .A (n_1490), .B (n_1492));
AOI22_X1 i_821 (.ZN (n_1492), .A1 (n_1308), .A2 (n_1491), .B1 (n_1307), .B2 (n_1304));
INV_X1 i_820 (.ZN (n_1491), .A (n_1309));
XNOR2_X1 i_819 (.ZN (n_1490), .A (n_1473), .B (n_1489));
XNOR2_X1 i_818 (.ZN (n_1489), .A (n_1487), .B (n_1488));
AOI22_X1 i_817 (.ZN (n_1488), .A1 (n_1337), .A2 (n_1351), .B1 (n_1350), .B2 (n_1342));
XNOR2_X1 i_816 (.ZN (n_1487), .A (n_1475), .B (n_1486));
XNOR2_X1 i_815 (.ZN (n_1486), .A (n_1326), .B (n_1338));
AOI22_X1 i_814 (.ZN (n_1475), .A1 (n_1144), .A2 (n_1474), .B1 (n_1196), .B2 (n_1145));
INV_X1 i_813 (.ZN (n_1474), .A (n_1288));
AOI22_X1 i_812 (.ZN (n_1473), .A1 (n_1380), .A2 (n_1391), .B1 (n_1472), .B2 (n_1379));
INV_X1 i_811 (.ZN (n_1472), .A (n_1356));
XNOR2_X1 i_810 (.ZN (n_1471), .A (n_1468), .B (n_1470));
AOI22_X1 i_809 (.ZN (n_1470), .A1 (n_1354), .A2 (n_1392), .B1 (n_1469), .B2 (n_1353));
INV_X1 i_808 (.ZN (n_1469), .A (n_1314));
XOR2_X1 i_807 (.Z (n_1468), .A (n_1430), .B (n_1467));
OAI21_X1 i_806 (.ZN (n_1467), .A (n_1466), .B1 (n_1431), .B2 (n_1465));
NAND2_X1 i_805 (.ZN (n_1466), .A1 (n_1431), .A2 (n_1465));
XOR2_X1 i_804 (.Z (n_1465), .A (n_1446), .B (n_1464));
XNOR2_X1 i_803 (.ZN (n_1464), .A (n_1458), .B (n_1463));
XNOR2_X1 i_802 (.ZN (n_1463), .A (n_1522), .B (n_1462));
NAND2_X1 i_801 (.ZN (n_1462), .A1 (A[8]), .A2 (B[17]));
XOR2_X1 i_800 (.Z (n_1458), .A (n_1451), .B (n_1457));
XNOR2_X1 i_799 (.ZN (n_1457), .A (n_1505), .B (n_1504));
XNOR2_X1 i_798 (.ZN (n_1451), .A (n_1371), .B (n_1372));
XNOR2_X1 i_797 (.ZN (n_1446), .A (n_1440), .B (n_1445));
XOR2_X1 i_796 (.Z (n_1445), .A (n_1526), .B (n_1341));
XNOR2_X1 i_795 (.ZN (n_1440), .A (n_1435), .B (n_1439));
XOR2_X1 i_794 (.Z (n_1439), .A (n_1437), .B (n_1438));
NAND2_X1 i_793 (.ZN (n_1438), .A1 (B[11]), .A2 (A[14]));
XNOR2_X1 i_792 (.ZN (n_1437), .A (n_1344), .B (n_1631));
XOR2_X1 i_791 (.Z (n_1435), .A (n_1433), .B (n_1434));
NAND2_X1 i_790 (.ZN (n_1434), .A1 (B[8]), .A2 (A[17]));
XNOR2_X1 i_789 (.ZN (n_1433), .A (n_1375), .B (n_1432));
NAND2_X1 i_788 (.ZN (n_1432), .A1 (B[6]), .A2 (A[19]));
AOI22_X1 i_787 (.ZN (n_1431), .A1 (n_1386), .A2 (n_1390), .B1 (n_1389), .B2 (n_1388));
XOR2_X1 i_786 (.Z (n_1430), .A (n_1428), .B (n_1429));
AOI22_X1 i_785 (.ZN (n_1429), .A1 (n_1336), .A2 (n_1352), .B1 (n_1316), .B2 (n_1335));
XOR2_X1 i_784 (.Z (n_1428), .A (n_1417), .B (n_1427));
XOR2_X1 i_783 (.Z (n_1427), .A (n_1423), .B (n_1442));
XOR2_X1 i_782 (.Z (n_1417), .A (n_1408), .B (n_1416));
XNOR2_X1 i_781 (.ZN (n_1416), .A (n_1501), .B (n_1461));
XNOR2_X1 i_780 (.ZN (n_1408), .A (n_1401), .B (n_1407));
XNOR2_X1 i_779 (.ZN (n_1407), .A (n_1362), .B (n_1365));
AOI22_X1 i_778 (.ZN (n_1401), .A1 (n_1236), .A2 (n_1385), .B1 (n_1263), .B2 (n_1400));
INV_X1 i_777 (.ZN (n_1400), .A (n_1239));
OAI21_X1 i_776 (.ZN (n_1399), .A (n_1284), .B1 (n_1398), .B2 (n_1285));
XNOR2_X1 i_775 (.ZN (Out[24]), .A (n_1287), .B (n_1398));
AOI21_X1 i_774 (.ZN (n_1398), .A (n_1397), .B1 (n_1396), .B2 (n_1394));
NOR2_X1 i_773 (.ZN (n_1397), .A1 (n_1394), .A2 (n_1396));
INV_X1 i_772 (.ZN (n_1396), .A (n_1395));
AOI22_X1 i_771 (.ZN (n_1395), .A1 (n_1278), .A2 (n_1246), .B1 (n_1247), .B2 (n_1277));
XOR2_X1 i_770 (.Z (n_1394), .A (n_1313), .B (n_1393));
XNOR2_X1 i_769 (.ZN (n_1393), .A (n_1354), .B (n_1392));
XOR2_X1 i_768 (.Z (n_1392), .A (n_1380), .B (n_1391));
XOR2_X1 i_767 (.Z (n_1391), .A (n_1386), .B (n_1390));
XOR2_X1 i_766 (.Z (n_1390), .A (n_1388), .B (n_1389));
AOI22_X1 i_765 (.ZN (n_1389), .A1 (n_1234), .A2 (n_1240), .B1 (n_1229), .B2 (n_1233));
OAI22_X1 i_764 (.ZN (n_1388), .A1 (n_1219), .A2 (n_1223), .B1 (n_1216), .B2 (n_1387));
INV_X1 i_763 (.ZN (n_1387), .A (n_1218));
XNOR2_X1 i_762 (.ZN (n_1386), .A (n_1236), .B (n_1385));
AOI22_X1 i_761 (.ZN (n_1385), .A1 (n_1270), .A2 (n_1267), .B1 (n_1268), .B2 (n_1269));
XNOR2_X1 i_760 (.ZN (n_1380), .A (n_1356), .B (n_1379));
OAI21_X1 i_759 (.ZN (n_1379), .A (n_1441), .B1 (n_1426), .B2 (n_1436));
AOI22_X1 i_758 (.ZN (n_1356), .A1 (n_1251), .A2 (n_1257), .B1 (n_1355), .B2 (n_1248));
INV_X1 i_757 (.ZN (n_1355), .A (n_1250));
XNOR2_X1 i_756 (.ZN (n_1354), .A (n_1314), .B (n_1353));
XOR2_X1 i_755 (.Z (n_1353), .A (n_1336), .B (n_1352));
XOR2_X1 i_754 (.Z (n_1352), .A (n_1337), .B (n_1351));
XOR2_X1 i_753 (.Z (n_1351), .A (n_1342), .B (n_1350));
XNOR2_X1 i_752 (.ZN (n_1350), .A (n_1347), .B (n_1482));
NAND2_X1 i_751 (.ZN (n_1347), .A1 (n_1484), .A2 (n_1485));
XNOR2_X1 i_750 (.ZN (n_1342), .A (n_1340), .B (n_1478));
NAND2_X1 i_749 (.ZN (n_1340), .A1 (n_1479), .A2 (n_1481));
AOI22_X1 i_748 (.ZN (n_1337), .A1 (n_1255), .A2 (n_1256), .B1 (n_1253), .B2 (n_1254));
XOR2_X1 i_747 (.Z (n_1336), .A (n_1316), .B (n_1335));
XOR2_X1 i_746 (.Z (n_1335), .A (n_1418), .B (n_1420));
AOI22_X1 i_745 (.ZN (n_1316), .A1 (n_1272), .A2 (n_1315), .B1 (n_1271), .B2 (n_1265));
INV_X1 i_744 (.ZN (n_1315), .A (n_1273));
AOI22_X1 i_743 (.ZN (n_1314), .A1 (n_1276), .A2 (n_1275), .B1 (n_1258), .B2 (n_1274));
XOR2_X1 i_742 (.Z (n_1313), .A (n_1310), .B (n_1312));
AOI22_X1 i_741 (.ZN (n_1312), .A1 (n_1244), .A2 (n_1311), .B1 (n_1210), .B2 (n_1243));
INV_X1 i_740 (.ZN (n_1311), .A (n_1245));
XOR2_X1 i_739 (.Z (n_1310), .A (n_1308), .B (n_1309));
AOI22_X1 i_738 (.ZN (n_1309), .A1 (n_1211), .A2 (n_1242), .B1 (n_1241), .B2 (n_1224));
XOR2_X1 i_737 (.Z (n_1308), .A (n_1304), .B (n_1307));
AOI22_X1 i_736 (.ZN (n_1307), .A1 (n_1208), .A2 (n_1030), .B1 (n_1306), .B2 (n_1207));
INV_X1 i_735 (.ZN (n_1306), .A (n_1189));
XOR2_X1 i_734 (.Z (n_1304), .A (n_1288), .B (n_1144));
AOI22_X1 i_733 (.ZN (n_1288), .A1 (n_1202), .A2 (n_1206), .B1 (n_1201), .B2 (n_1195));
NAND2_X1 i_732 (.ZN (n_1287), .A1 (n_1284), .A2 (n_1286));
INV_X1 i_731 (.ZN (n_1286), .A (n_1285));
NOR4_X1 i_730 (.ZN (n_1285), .A1 (n_1090), .A2 (n_1185), .A3 (n_1283), .A4 (n_1279));
OAI21_X1 i_729 (.ZN (n_1284), .A (n_1282), .B1 (n_1283), .B2 (n_1279));
INV_X1 i_728 (.ZN (n_1283), .A (n_1188));
OAI21_X1 i_727 (.ZN (n_1282), .A (n_1280), .B1 (n_1187), .B2 (n_1281));
XNOR2_X1 i_726 (.ZN (Out[23]), .A (n_1187), .B (n_1281));
XOR2_X1 i_725 (.Z (n_1281), .A (n_1280), .B (n_1185));
XNOR2_X1 i_724 (.ZN (n_1280), .A (n_1188), .B (n_1279));
XOR2_X1 i_723 (.Z (n_1279), .A (n_1246), .B (n_1278));
XOR2_X1 i_722 (.Z (n_1278), .A (n_1247), .B (n_1277));
XNOR2_X1 i_721 (.ZN (n_1277), .A (n_1275), .B (n_1276));
AOI22_X1 i_720 (.ZN (n_1276), .A1 (n_1142), .A2 (n_1178), .B1 (n_1163), .B2 (n_1177));
XOR2_X1 i_719 (.Z (n_1275), .A (n_1258), .B (n_1274));
XOR2_X1 i_718 (.Z (n_1274), .A (n_1272), .B (n_1273));
AOI22_X1 i_717 (.ZN (n_1273), .A1 (n_1172), .A2 (n_1176), .B1 (n_1171), .B2 (n_1167));
XOR2_X1 i_716 (.Z (n_1272), .A (n_1265), .B (n_1271));
XNOR2_X1 i_715 (.ZN (n_1271), .A (n_1267), .B (n_1270));
XOR2_X1 i_714 (.Z (n_1270), .A (n_1268), .B (n_1269));
OAI22_X1 i_713 (.ZN (n_1269), .A1 (n_1165), .A2 (n_1166), .B1 (n_1051), .B2 (n_1231));
OAI22_X1 i_712 (.ZN (n_1268), .A1 (n_1169), .A2 (n_1170), .B1 (n_1060), .B2 (n_1168));
OAI33_X1 i_711 (.ZN (n_1267), .A1 (n_1174), .A2 (n_99), .A3 (n_1711), .B1 (n_1209)
    , .B2 (n_423), .B3 (n_1232));
XOR2_X1 i_710 (.Z (n_1265), .A (n_1292), .B (n_1264));
XOR2_X1 i_709 (.Z (n_1258), .A (n_1251), .B (n_1257));
XNOR2_X1 i_708 (.ZN (n_1257), .A (n_1255), .B (n_1256));
AOI22_X1 i_707 (.ZN (n_1256), .A1 (n_1061), .A2 (n_1056), .B1 (n_1063), .B2 (n_1062));
XOR2_X1 i_706 (.Z (n_1255), .A (n_1253), .B (n_1254));
AND2_X1 i_705 (.ZN (n_1254), .A1 (n_1134), .A2 (n_1130));
AOI22_X1 i_704 (.ZN (n_1253), .A1 (n_1139), .A2 (n_1140), .B1 (n_1252), .B2 (n_1138));
INV_X1 i_703 (.ZN (n_1252), .A (n_1137));
XNOR2_X1 i_702 (.ZN (n_1251), .A (n_1248), .B (n_1250));
AOI22_X1 i_701 (.ZN (n_1250), .A1 (n_955), .A2 (n_945), .B1 (n_1249), .B2 (n_978));
INV_X1 i_700 (.ZN (n_1249), .A (n_999));
AOI22_X1 i_699 (.ZN (n_1248), .A1 (n_1156), .A2 (n_1162), .B1 (n_1149), .B2 (n_1155));
AOI22_X1 i_698 (.ZN (n_1247), .A1 (n_1180), .A2 (n_1181), .B1 (n_1179), .B2 (n_1124));
XOR2_X1 i_697 (.Z (n_1246), .A (n_1244), .B (n_1245));
AOI22_X1 i_696 (.ZN (n_1245), .A1 (n_1094), .A2 (n_1107), .B1 (n_1106), .B2 (n_1105));
XOR2_X1 i_695 (.Z (n_1244), .A (n_1210), .B (n_1243));
XOR2_X1 i_694 (.Z (n_1243), .A (n_1211), .B (n_1242));
XOR2_X1 i_693 (.Z (n_1242), .A (n_1224), .B (n_1241));
XNOR2_X1 i_692 (.ZN (n_1241), .A (n_1234), .B (n_1240));
XNOR2_X1 i_691 (.ZN (n_1240), .A (n_1238), .B (n_1214));
NAND2_X1 i_690 (.ZN (n_1238), .A1 (n_1220), .A2 (n_1237));
INV_X1 i_689 (.ZN (n_1237), .A (n_1221));
XOR2_X1 i_688 (.Z (n_1234), .A (n_1229), .B (n_1233));
XNOR2_X1 i_687 (.ZN (n_1233), .A (n_1150), .B (n_1148));
XOR2_X1 i_686 (.Z (n_1229), .A (n_1158), .B (n_1157));
XOR2_X1 i_685 (.Z (n_1224), .A (n_1219), .B (n_1223));
XNOR2_X1 i_684 (.ZN (n_1223), .A (n_1192), .B (n_1191));
XOR2_X1 i_683 (.Z (n_1219), .A (n_1216), .B (n_1218));
AOI21_X1 i_682 (.ZN (n_1218), .A (n_947), .B1 (n_950), .B2 (n_1217));
INV_X1 i_681 (.ZN (n_1217), .A (n_948));
XOR2_X1 i_680 (.Z (n_1216), .A (n_1215), .B (n_949));
NOR2_X1 i_679 (.ZN (n_1215), .A1 (n_1329), .A2 (n_1327));
AOI22_X1 i_678 (.ZN (n_1211), .A1 (n_903), .A2 (n_1123), .B1 (n_904), .B2 (n_944));
XOR2_X1 i_677 (.Z (n_1210), .A (n_1208), .B (n_1031));
XNOR2_X1 i_676 (.ZN (n_1208), .A (n_1189), .B (n_1207));
XOR2_X1 i_675 (.Z (n_1207), .A (n_1202), .B (n_1206));
XNOR2_X1 i_674 (.ZN (n_1206), .A (n_1260), .B (n_1259));
XOR2_X1 i_673 (.Z (n_1202), .A (n_1195), .B (n_1201));
XNOR2_X1 i_672 (.ZN (n_1201), .A (n_1226), .B (n_1225));
XNOR2_X1 i_671 (.ZN (n_1195), .A (n_1200), .B (n_1199));
AOI22_X1 i_670 (.ZN (n_1189), .A1 (n_1136), .A2 (n_1141), .B1 (n_1126), .B2 (n_1135));
AOI22_X1 i_669 (.ZN (n_1188), .A1 (n_1109), .A2 (n_1182), .B1 (n_1093), .B2 (n_1108));
OAI21_X1 i_668 (.ZN (n_1187), .A (n_1090), .B1 (n_1088), .B2 (n_1186));
XOR2_X1 i_667 (.Z (Out[22]), .A (n_1091), .B (n_1186));
OAI21_X1 i_666 (.ZN (n_1186), .A (n_1185), .B1 (n_1184), .B2 (n_1183));
NAND2_X1 i_665 (.ZN (n_1185), .A1 (n_1183), .A2 (n_1184));
OAI22_X1 i_664 (.ZN (n_1184), .A1 (n_1043), .A2 (n_1076), .B1 (n_1045), .B2 (n_1075));
XNOR2_X1 i_663 (.ZN (n_1183), .A (n_1109), .B (n_1182));
XNOR2_X1 i_662 (.ZN (n_1182), .A (n_1180), .B (n_1181));
AOI22_X1 i_661 (.ZN (n_1181), .A1 (n_1067), .A2 (n_1074), .B1 (n_1047), .B2 (n_1066));
XOR2_X1 i_660 (.Z (n_1180), .A (n_1124), .B (n_1179));
XNOR2_X1 i_659 (.ZN (n_1179), .A (n_1142), .B (n_1178));
XOR2_X1 i_658 (.Z (n_1178), .A (n_1163), .B (n_1177));
XOR2_X1 i_657 (.Z (n_1177), .A (n_1172), .B (n_1176));
XNOR2_X1 i_656 (.ZN (n_1176), .A (n_1174), .B (n_1175));
NAND2_X1 i_655 (.ZN (n_1175), .A1 (A[3]), .A2 (B[19]));
XNOR2_X1 i_654 (.ZN (n_1174), .A (n_889), .B (n_1209));
XOR2_X1 i_653 (.Z (n_1172), .A (n_1167), .B (n_1171));
XNOR2_X1 i_652 (.ZN (n_1171), .A (n_1169), .B (n_1170));
NAND2_X1 i_651 (.ZN (n_1170), .A1 (A[9]), .A2 (B[13]));
XNOR2_X1 i_650 (.ZN (n_1169), .A (n_1060), .B (n_1168));
NAND2_X1 i_649 (.ZN (n_1168), .A1 (B[11]), .A2 (A[11]));
XNOR2_X1 i_648 (.ZN (n_1167), .A (n_1165), .B (n_1166));
NAND2_X1 i_647 (.ZN (n_1166), .A1 (A[6]), .A2 (B[16]));
XNOR2_X1 i_646 (.ZN (n_1165), .A (n_1051), .B (n_1231));
XOR2_X1 i_645 (.Z (n_1163), .A (n_1156), .B (n_1162));
XOR2_X1 i_644 (.Z (n_1162), .A (n_1289), .B (n_1173));
XOR2_X1 i_643 (.Z (n_1156), .A (n_1149), .B (n_1155));
XNOR2_X1 i_642 (.ZN (n_1155), .A (n_1296), .B (n_1295));
XNOR2_X1 i_641 (.ZN (n_1149), .A (n_1301), .B (n_1300));
XOR2_X1 i_640 (.Z (n_1142), .A (n_1136), .B (n_1141));
XNOR2_X1 i_639 (.ZN (n_1141), .A (n_1139), .B (n_1140));
AOI21_X1 i_638 (.ZN (n_1140), .A (n_896), .B1 (n_902), .B2 (n_888));
XNOR2_X1 i_637 (.ZN (n_1139), .A (n_1137), .B (n_1138));
AOI21_X1 i_636 (.ZN (n_1138), .A (n_884), .B1 (n_860), .B2 (n_855));
AOI21_X1 i_635 (.ZN (n_1137), .A (n_1050), .B1 (n_1048), .B2 (n_1036));
XOR2_X1 i_634 (.Z (n_1136), .A (n_1126), .B (n_1135));
NAND2_X1 i_633 (.ZN (n_1135), .A1 (n_1133), .A2 (n_1134));
OR3_X1 i_632 (.ZN (n_1134), .A1 (n_1131), .A2 (n_1132), .A3 (n_1127));
OAI21_X1 i_631 (.ZN (n_1133), .A (n_1127), .B1 (n_1131), .B2 (n_1132));
AOI22_X1 i_630 (.ZN (n_1132), .A1 (A[1]), .A2 (B[21]), .B1 (A[2]), .B2 (B[20]));
INV_X1 i_629 (.ZN (n_1131), .A (n_1130));
NAND3_X1 i_628 (.ZN (n_1130), .A1 (n_1530), .A2 (A[1]), .A3 (B[20]));
NAND2_X1 i_627 (.ZN (n_1127), .A1 (A[0]), .A2 (B[22]));
AOI22_X1 i_626 (.ZN (n_1126), .A1 (n_980), .A2 (n_1125), .B1 (n_979), .B2 (n_977));
INV_X1 i_625 (.ZN (n_1125), .A (n_982));
XNOR2_X1 i_624 (.ZN (n_1124), .A (n_903), .B (n_1123));
AOI22_X1 i_623 (.ZN (n_1123), .A1 (n_983), .A2 (n_901), .B1 (n_887), .B2 (n_899));
XOR2_X1 i_622 (.Z (n_1109), .A (n_1093), .B (n_1108));
XNOR2_X1 i_621 (.ZN (n_1108), .A (n_1094), .B (n_1107));
XOR2_X1 i_620 (.Z (n_1107), .A (n_1105), .B (n_1106));
OAI21_X1 i_619 (.ZN (n_1106), .A (n_1071), .B1 (n_1072), .B2 (n_1073));
XNOR2_X1 i_618 (.ZN (n_1105), .A (n_1032), .B (n_1096));
AOI22_X1 i_617 (.ZN (n_1094), .A1 (n_1020), .A2 (n_1037), .B1 (n_997), .B2 (n_1019));
AOI22_X1 i_616 (.ZN (n_1093), .A1 (n_1041), .A2 (n_1042), .B1 (n_1038), .B2 (n_1092));
INV_X1 i_615 (.ZN (n_1092), .A (n_1040));
NAND2_X1 i_614 (.ZN (n_1091), .A1 (n_1089), .A2 (n_1090));
NAND2_X1 i_613 (.ZN (n_1090), .A1 (n_1086), .A2 (n_1087));
INV_X1 i_612 (.ZN (n_1089), .A (n_1088));
NOR2_X1 i_611 (.ZN (n_1088), .A1 (n_1086), .A2 (n_1087));
INV_X1 i_610 (.ZN (n_1087), .A (n_1079));
OAI21_X1 i_609 (.ZN (n_1086), .A (n_1085), .B1 (n_975), .B2 (n_1082));
INV_X1 i_608 (.ZN (n_1085), .A (n_1083));
XNOR2_X1 i_607 (.ZN (Out[21]), .A (n_975), .B (n_1084));
NOR2_X1 i_606 (.ZN (n_1084), .A1 (n_1082), .A2 (n_1083));
NOR2_X1 i_605 (.ZN (n_1083), .A1 (n_1080), .A2 (n_1081));
AND2_X1 i_604 (.ZN (n_1082), .A1 (n_1080), .A2 (n_1081));
INV_X1 i_603 (.ZN (n_1081), .A (n_973));
OAI21_X1 i_602 (.ZN (n_1080), .A (n_1079), .B1 (n_1077), .B2 (n_1078));
NAND2_X1 i_601 (.ZN (n_1079), .A1 (n_1077), .A2 (n_1078));
OAI21_X1 i_600 (.ZN (n_1078), .A (n_935), .B1 (n_936), .B2 (n_965));
XOR2_X1 i_599 (.Z (n_1077), .A (n_1043), .B (n_1076));
XNOR2_X1 i_598 (.ZN (n_1076), .A (n_1045), .B (n_1075));
XOR2_X1 i_597 (.Z (n_1075), .A (n_1067), .B (n_1074));
XNOR2_X1 i_596 (.ZN (n_1074), .A (n_1072), .B (n_1073));
AOI22_X1 i_595 (.ZN (n_1073), .A1 (n_923), .A2 (n_930), .B1 (n_917), .B2 (n_922));
OAI21_X1 i_594 (.ZN (n_1072), .A (n_1071), .B1 (n_1069), .B2 (n_1070));
NAND2_X1 i_593 (.ZN (n_1071), .A1 (n_1069), .A2 (n_1070));
AOI22_X1 i_592 (.ZN (n_1070), .A1 (n_908), .A2 (n_914), .B1 (n_907), .B2 (n_900));
AOI22_X1 i_591 (.ZN (n_1069), .A1 (n_883), .A2 (n_890), .B1 (n_881), .B2 (n_1068));
INV_X1 i_590 (.ZN (n_1068), .A (n_882));
XOR2_X1 i_589 (.Z (n_1067), .A (n_1047), .B (n_1066));
XNOR2_X1 i_588 (.ZN (n_1066), .A (n_940), .B (n_905));
AOI22_X1 i_587 (.ZN (n_1047), .A1 (n_891), .A2 (n_894), .B1 (n_1046), .B2 (n_893));
INV_X1 i_586 (.ZN (n_1046), .A (n_892));
OAI22_X1 i_585 (.ZN (n_1045), .A1 (n_959), .A2 (n_964), .B1 (n_1044), .B2 (n_963));
INV_X1 i_584 (.ZN (n_1044), .A (n_960));
XNOR2_X1 i_583 (.ZN (n_1043), .A (n_1041), .B (n_1042));
AOI22_X1 i_582 (.ZN (n_1042), .A1 (n_916), .A2 (n_931), .B1 (n_895), .B2 (n_915));
XNOR2_X1 i_581 (.ZN (n_1041), .A (n_1038), .B (n_1040));
AOI22_X1 i_580 (.ZN (n_1040), .A1 (n_957), .A2 (n_958), .B1 (n_1039), .B2 (n_956));
INV_X1 i_579 (.ZN (n_1039), .A (n_937));
XNOR2_X1 i_578 (.ZN (n_1038), .A (n_1020), .B (n_1037));
XNOR2_X1 i_577 (.ZN (n_1037), .A (n_1103), .B (n_1097));
XOR2_X1 i_576 (.Z (n_1020), .A (n_997), .B (n_1019));
XOR2_X1 i_575 (.Z (n_1019), .A (n_1012), .B (n_1035));
NAND2_X1 i_574 (.ZN (n_1012), .A1 (n_1010), .A2 (n_1053));
INV_X1 i_573 (.ZN (n_1010), .A (n_1052));
XNOR2_X1 i_572 (.ZN (n_997), .A (n_983), .B (n_901));
XNOR2_X1 i_571 (.ZN (n_983), .A (n_980), .B (n_982));
AOI22_X1 i_570 (.ZN (n_982), .A1 (n_920), .A2 (n_921), .B1 (n_918), .B2 (n_981));
INV_X1 i_569 (.ZN (n_981), .A (n_919));
XOR2_X1 i_568 (.Z (n_980), .A (n_977), .B (n_979));
OAI33_X1 i_567 (.ZN (n_979), .A1 (n_928), .A2 (n_99), .A3 (n_1232), .B1 (n_939), .B2 (n_423), .B3 (n_560));
NAND2_X1 i_566 (.ZN (n_977), .A1 (n_909), .A2 (n_976));
INV_X1 i_565 (.ZN (n_976), .A (n_912));
AOI21_X1 i_564 (.ZN (n_975), .A (n_967), .B1 (n_974), .B2 (n_969));
XNOR2_X1 i_563 (.ZN (Out[20]), .A (n_970), .B (n_974));
AOI21_X1 i_562 (.ZN (n_974), .A (n_973), .B1 (n_874), .B2 (n_972));
NOR2_X1 i_561 (.ZN (n_973), .A1 (n_874), .A2 (n_972));
OAI22_X1 i_560 (.ZN (n_972), .A1 (n_870), .A2 (n_971), .B1 (n_828), .B2 (n_869));
INV_X1 i_559 (.ZN (n_971), .A (n_871));
NAND2_X1 i_558 (.ZN (n_970), .A1 (n_968), .A2 (n_969));
NAND2_X1 i_557 (.ZN (n_969), .A1 (n_878), .A2 (n_966));
INV_X1 i_556 (.ZN (n_968), .A (n_967));
NOR2_X1 i_555 (.ZN (n_967), .A1 (n_878), .A2 (n_966));
XNOR2_X1 i_554 (.ZN (n_966), .A (n_936), .B (n_965));
XOR2_X1 i_553 (.Z (n_965), .A (n_959), .B (n_964));
XOR2_X1 i_552 (.Z (n_964), .A (n_960), .B (n_963));
AOI22_X1 i_551 (.ZN (n_963), .A1 (n_796), .A2 (n_811), .B1 (n_961), .B2 (n_962));
INV_X1 i_550 (.ZN (n_962), .A (n_795));
INV_X1 i_549 (.ZN (n_961), .A (n_794));
OAI21_X1 i_548 (.ZN (n_960), .A (n_867), .B1 (n_832), .B2 (n_868));
XOR2_X1 i_547 (.Z (n_959), .A (n_957), .B (n_958));
AOI22_X1 i_546 (.ZN (n_958), .A1 (n_801), .A2 (n_810), .B1 (n_809), .B2 (n_805));
XNOR2_X1 i_545 (.ZN (n_957), .A (n_937), .B (n_956));
XNOR2_X1 i_544 (.ZN (n_956), .A (n_924), .B (n_906));
AOI22_X1 i_543 (.ZN (n_937), .A1 (n_820), .A2 (n_822), .B1 (n_819), .B2 (n_813));
OAI21_X1 i_542 (.ZN (n_936), .A (n_935), .B1 (n_932), .B2 (n_934));
NAND2_X1 i_541 (.ZN (n_935), .A1 (n_932), .A2 (n_934));
OAI21_X1 i_540 (.ZN (n_934), .A (n_824), .B1 (n_933), .B2 (n_827));
INV_X1 i_539 (.ZN (n_933), .A (n_825));
XNOR2_X1 i_538 (.ZN (n_932), .A (n_916), .B (n_931));
XNOR2_X1 i_537 (.ZN (n_931), .A (n_923), .B (n_930));
XOR2_X1 i_536 (.Z (n_930), .A (n_1117), .B (n_1113));
XOR2_X1 i_535 (.Z (n_923), .A (n_917), .B (n_922));
XOR2_X1 i_534 (.Z (n_922), .A (n_920), .B (n_921));
OAI22_X1 i_533 (.ZN (n_921), .A1 (n_807), .A2 (n_808), .B1 (n_716), .B2 (n_806));
XNOR2_X1 i_532 (.ZN (n_920), .A (n_918), .B (n_919));
AOI21_X1 i_531 (.ZN (n_919), .A (n_861), .B1 (n_863), .B2 (n_864));
OAI22_X1 i_530 (.ZN (n_918), .A1 (n_804), .A2 (n_722), .B1 (n_913), .B2 (n_803));
OAI22_X1 i_529 (.ZN (n_917), .A1 (n_797), .A2 (n_800), .B1 (n_798), .B2 (n_799));
XOR2_X1 i_528 (.Z (n_916), .A (n_895), .B (n_915));
XOR2_X1 i_527 (.Z (n_915), .A (n_908), .B (n_914));
XOR2_X1 i_526 (.Z (n_914), .A (n_1022), .B (n_1021));
XOR2_X1 i_525 (.Z (n_908), .A (n_900), .B (n_907));
XNOR2_X1 i_524 (.ZN (n_907), .A (n_995), .B (n_994));
XOR2_X1 i_523 (.Z (n_900), .A (n_1013), .B (n_1011));
XNOR2_X1 i_522 (.ZN (n_895), .A (n_891), .B (n_894));
XNOR2_X1 i_521 (.ZN (n_894), .A (n_892), .B (n_893));
AOI22_X1 i_520 (.ZN (n_893), .A1 (n_859), .A2 (n_865), .B1 (n_854), .B2 (n_858));
AOI22_X1 i_519 (.ZN (n_892), .A1 (n_840), .A2 (n_834), .B1 (n_847), .B2 (n_841));
XNOR2_X1 i_518 (.ZN (n_891), .A (n_883), .B (n_890));
XNOR2_X1 i_517 (.ZN (n_890), .A (n_990), .B (n_989));
XNOR2_X1 i_516 (.ZN (n_883), .A (n_881), .B (n_882));
AOI21_X1 i_515 (.ZN (n_882), .A (n_843), .B1 (n_846), .B2 (n_844));
AOI22_X1 i_514 (.ZN (n_881), .A1 (n_818), .A2 (n_816), .B1 (n_815), .B2 (n_814));
OAI21_X1 i_513 (.ZN (Out[19]), .A (n_879), .B1 (n_875), .B2 (n_880));
INV_X1 i_512 (.ZN (n_880), .A (n_877));
OAI21_X1 i_511 (.ZN (n_879), .A (n_878), .B1 (n_792), .B2 (n_876));
OAI21_X1 i_510 (.ZN (n_878), .A (n_792), .B1 (n_876), .B2 (n_877));
NOR2_X1 i_509 (.ZN (n_877), .A1 (n_710), .A2 (n_790));
INV_X1 i_508 (.ZN (n_876), .A (n_875));
OAI21_X1 i_507 (.ZN (n_875), .A (n_874), .B1 (n_872), .B2 (n_873));
NAND2_X1 i_506 (.ZN (n_874), .A1 (n_872), .A2 (n_873));
AOI22_X1 i_505 (.ZN (n_873), .A1 (n_786), .A2 (n_753), .B1 (n_712), .B2 (n_752));
XOR2_X1 i_504 (.Z (n_872), .A (n_870), .B (n_871));
AOI22_X1 i_503 (.ZN (n_871), .A1 (n_768), .A2 (n_785), .B1 (n_754), .B2 (n_767));
XNOR2_X1 i_502 (.ZN (n_870), .A (n_828), .B (n_869));
XNOR2_X1 i_501 (.ZN (n_869), .A (n_832), .B (n_868));
OAI21_X1 i_500 (.ZN (n_868), .A (n_867), .B1 (n_866), .B2 (n_833));
NAND2_X1 i_499 (.ZN (n_867), .A1 (n_833), .A2 (n_866));
XOR2_X1 i_498 (.Z (n_866), .A (n_859), .B (n_865));
XNOR2_X1 i_497 (.ZN (n_865), .A (n_863), .B (n_864));
NOR2_X1 i_496 (.ZN (n_864), .A1 (n_170), .A2 (n_229));
NOR2_X1 i_495 (.ZN (n_863), .A1 (n_861), .A2 (n_862));
AOI22_X1 i_494 (.ZN (n_862), .A1 (A[7]), .A2 (B[12]), .B1 (A[8]), .B2 (B[11]));
NOR2_X1 i_493 (.ZN (n_861), .A1 (n_743), .A2 (n_1008));
XOR2_X1 i_492 (.Z (n_859), .A (n_854), .B (n_858));
XNOR2_X1 i_491 (.ZN (n_858), .A (n_1115), .B (n_1114));
XOR2_X1 i_490 (.Z (n_854), .A (n_1120), .B (n_1017));
XOR2_X1 i_489 (.Z (n_828), .A (n_826), .B (n_827));
OAI21_X1 i_488 (.ZN (n_827), .A (n_748), .B1 (n_751), .B2 (n_749));
NAND2_X1 i_487 (.ZN (n_826), .A1 (n_824), .A2 (n_825));
NAND2_X1 i_486 (.ZN (n_825), .A1 (n_812), .A2 (n_823));
OR2_X1 i_485 (.ZN (n_824), .A1 (n_812), .A2 (n_823));
XNOR2_X1 i_484 (.ZN (n_823), .A (n_820), .B (n_822));
OAI22_X1 i_483 (.ZN (n_822), .A1 (n_694), .A2 (n_761), .B1 (n_760), .B2 (n_821));
INV_X1 i_482 (.ZN (n_821), .A (n_750));
XOR2_X1 i_481 (.Z (n_820), .A (n_813), .B (n_819));
XOR2_X1 i_480 (.Z (n_819), .A (n_816), .B (n_818));
OAI33_X1 i_479 (.ZN (n_818), .A1 (n_744), .A2 (n_170), .A3 (n_1676), .B1 (n_743), .B2 (n_2243), .B3 (n_458));
XOR2_X1 i_478 (.Z (n_816), .A (n_814), .B (n_815));
OAI22_X1 i_477 (.ZN (n_815), .A1 (n_739), .A2 (n_740), .B1 (n_1128), .B2 (n_738));
OAI21_X1 i_476 (.ZN (n_814), .A (n_732), .B1 (n_734), .B2 (n_735));
AOI22_X1 i_475 (.ZN (n_813), .A1 (n_742), .A2 (n_746), .B1 (n_736), .B2 (n_741));
XOR2_X1 i_474 (.Z (n_812), .A (n_796), .B (n_811));
XOR2_X1 i_473 (.Z (n_811), .A (n_801), .B (n_810));
XOR2_X1 i_472 (.Z (n_810), .A (n_805), .B (n_809));
XNOR2_X1 i_471 (.ZN (n_809), .A (n_807), .B (n_808));
NAND2_X1 i_470 (.ZN (n_808), .A1 (A[3]), .A2 (B[16]));
XNOR2_X1 i_469 (.ZN (n_807), .A (n_716), .B (n_806));
NAND2_X1 i_468 (.ZN (n_806), .A1 (A[4]), .A2 (B[15]));
XNOR2_X1 i_467 (.ZN (n_805), .A (n_804), .B (n_722));
XNOR2_X1 i_466 (.ZN (n_804), .A (n_913), .B (n_803));
NAND2_X1 i_465 (.ZN (n_803), .A1 (A[0]), .A2 (B[19]));
XNOR2_X1 i_464 (.ZN (n_801), .A (n_797), .B (n_800));
XNOR2_X1 i_463 (.ZN (n_800), .A (n_798), .B (n_799));
AOI21_X1 i_462 (.ZN (n_799), .A (n_723), .B1 (n_725), .B2 (n_727));
AOI21_X1 i_461 (.ZN (n_798), .A (n_717), .B1 (n_719), .B2 (n_720));
AOI22_X1 i_460 (.ZN (n_797), .A1 (n_757), .A2 (n_758), .B1 (n_756), .B2 (n_755));
XOR2_X1 i_459 (.Z (n_796), .A (n_794), .B (n_795));
AOI22_X1 i_458 (.ZN (n_795), .A1 (n_715), .A2 (n_729), .B1 (n_721), .B2 (n_728));
AOI22_X1 i_457 (.ZN (n_794), .A1 (n_765), .A2 (n_793), .B1 (n_764), .B2 (n_759));
INV_X1 i_456 (.ZN (n_793), .A (n_766));
OAI211_X1 i_455 (.ZN (n_792), .A (n_710), .B (n_790), .C1 (n_791), .C2 (n_789));
INV_X1 i_454 (.ZN (n_791), .A (n_709));
NAND2_X1 i_453 (.ZN (n_790), .A1 (n_787), .A2 (n_788));
XOR2_X1 i_452 (.Z (Out[18]), .A (n_711), .B (n_789));
XNOR2_X1 i_451 (.ZN (n_789), .A (n_787), .B (n_788));
OAI21_X1 i_450 (.ZN (n_788), .A (n_701), .B1 (n_635), .B2 (n_673));
XNOR2_X1 i_449 (.ZN (n_787), .A (n_753), .B (n_786));
XNOR2_X1 i_448 (.ZN (n_786), .A (n_768), .B (n_785));
XOR2_X1 i_447 (.Z (n_785), .A (n_802), .B (n_831));
XOR2_X1 i_446 (.Z (n_768), .A (n_754), .B (n_767));
XOR2_X1 i_445 (.Z (n_767), .A (n_765), .B (n_766));
AOI22_X1 i_444 (.ZN (n_766), .A1 (n_653), .A2 (n_657), .B1 (n_644), .B2 (n_652));
XOR2_X1 i_443 (.Z (n_765), .A (n_759), .B (n_764));
XNOR2_X1 i_442 (.ZN (n_764), .A (n_849), .B (n_848));
XNOR2_X1 i_441 (.ZN (n_759), .A (n_757), .B (n_758));
OAI22_X1 i_440 (.ZN (n_758), .A1 (n_655), .A2 (n_656), .B1 (n_599), .B2 (n_654));
XOR2_X1 i_439 (.Z (n_757), .A (n_755), .B (n_756));
OAI21_X1 i_438 (.ZN (n_756), .A (n_649), .B1 (n_650), .B2 (n_651));
OAI21_X1 i_437 (.ZN (n_755), .A (n_639), .B1 (n_642), .B2 (n_643));
AOI22_X1 i_436 (.ZN (n_754), .A1 (n_659), .A2 (n_672), .B1 (n_637), .B2 (n_658));
XOR2_X1 i_435 (.Z (n_753), .A (n_712), .B (n_752));
XOR2_X1 i_434 (.Z (n_752), .A (n_749), .B (n_751));
AOI22_X1 i_433 (.ZN (n_751), .A1 (n_611), .A2 (n_459), .B1 (n_606), .B2 (n_610));
OAI21_X1 i_432 (.ZN (n_749), .A (n_748), .B1 (n_730), .B2 (n_747));
NAND2_X1 i_431 (.ZN (n_748), .A1 (n_730), .A2 (n_747));
XOR2_X1 i_430 (.Z (n_747), .A (n_742), .B (n_746));
XNOR2_X1 i_429 (.ZN (n_746), .A (n_744), .B (n_745));
NAND2_X1 i_428 (.ZN (n_745), .A1 (A[6]), .A2 (B[12]));
XNOR2_X1 i_427 (.ZN (n_744), .A (n_638), .B (n_743));
NAND2_X1 i_426 (.ZN (n_743), .A1 (A[7]), .A2 (B[11]));
XOR2_X1 i_425 (.Z (n_742), .A (n_736), .B (n_741));
XNOR2_X1 i_424 (.ZN (n_741), .A (n_739), .B (n_740));
NAND2_X1 i_423 (.ZN (n_740), .A1 (B[6]), .A2 (A[12]));
XNOR2_X1 i_422 (.ZN (n_739), .A (n_1128), .B (n_738));
NAND2_X1 i_421 (.ZN (n_738), .A1 (B[4]), .A2 (A[14]));
XNOR2_X1 i_420 (.ZN (n_736), .A (n_734), .B (n_735));
NAND2_X1 i_419 (.ZN (n_735), .A1 (A[9]), .A2 (B[9]));
NAND2_X1 i_418 (.ZN (n_734), .A1 (n_732), .A2 (n_733));
OAI22_X1 i_417 (.ZN (n_733), .A1 (n_425), .A2 (n_1339), .B1 (n_1955), .B2 (n_1235));
OR3_X1 i_416 (.ZN (n_732), .A1 (n_1116), .A2 (n_1955), .A3 (n_1339));
XOR2_X1 i_415 (.Z (n_730), .A (n_715), .B (n_729));
XOR2_X1 i_414 (.Z (n_729), .A (n_721), .B (n_728));
XNOR2_X1 i_413 (.ZN (n_728), .A (n_725), .B (n_727));
NOR2_X1 i_412 (.ZN (n_727), .A1 (n_31), .A2 (n_1532));
NOR2_X1 i_411 (.ZN (n_725), .A1 (n_723), .A2 (n_724));
AOI22_X1 i_410 (.ZN (n_724), .A1 (A[1]), .A2 (B[17]), .B1 (A[2]), .B2 (B[16]));
NOR2_X1 i_409 (.ZN (n_723), .A1 (n_607), .A2 (n_722));
NAND2_X1 i_408 (.ZN (n_722), .A1 (A[2]), .A2 (B[17]));
XNOR2_X1 i_407 (.ZN (n_721), .A (n_719), .B (n_720));
NOR2_X1 i_406 (.ZN (n_720), .A1 (n_99), .A2 (n_560));
NOR2_X1 i_405 (.ZN (n_719), .A1 (n_717), .A2 (n_718));
AOI22_X1 i_404 (.ZN (n_718), .A1 (A[4]), .A2 (B[14]), .B1 (A[5]), .B2 (B[13]));
NOR2_X1 i_403 (.ZN (n_717), .A1 (n_654), .A2 (n_716));
NAND2_X1 i_402 (.ZN (n_716), .A1 (A[5]), .A2 (B[14]));
AOI22_X1 i_401 (.ZN (n_715), .A1 (n_713), .A2 (n_605), .B1 (n_714), .B2 (n_604));
INV_X1 i_400 (.ZN (n_714), .A (n_598));
INV_X1 i_399 (.ZN (n_713), .A (n_582));
AOI22_X1 i_398 (.ZN (n_712), .A1 (n_698), .A2 (n_699), .B1 (n_688), .B2 (n_697));
NAND2_X1 i_397 (.ZN (n_711), .A1 (n_709), .A2 (n_710));
OR2_X1 i_396 (.ZN (n_710), .A1 (n_708), .A2 (n_633));
NAND2_X1 i_395 (.ZN (n_709), .A1 (n_708), .A2 (n_633));
INV_X1 i_394 (.ZN (n_708), .A (n_707));
OAI21_X1 i_393 (.ZN (n_707), .A (n_703), .B1 (n_631), .B2 (n_706));
INV_X1 i_392 (.ZN (n_706), .A (n_704));
XOR2_X1 i_391 (.Z (Out[17]), .A (n_631), .B (n_705));
NAND2_X1 i_390 (.ZN (n_705), .A1 (n_703), .A2 (n_704));
NAND2_X1 i_389 (.ZN (n_704), .A1 (n_634), .A2 (n_702));
OR2_X1 i_388 (.ZN (n_703), .A1 (n_634), .A2 (n_702));
OAI21_X1 i_387 (.ZN (n_702), .A (n_701), .B1 (n_674), .B2 (n_700));
NAND2_X1 i_386 (.ZN (n_701), .A1 (n_674), .A2 (n_700));
XOR2_X1 i_385 (.Z (n_700), .A (n_698), .B (n_699));
AOI22_X1 i_384 (.ZN (n_699), .A1 (n_554), .A2 (n_585), .B1 (n_563), .B2 (n_584));
XOR2_X1 i_383 (.Z (n_698), .A (n_688), .B (n_697));
XNOR2_X1 i_382 (.ZN (n_697), .A (n_777), .B (n_783));
XOR2_X1 i_381 (.Z (n_688), .A (n_611), .B (n_460));
XOR2_X1 i_380 (.Z (n_674), .A (n_635), .B (n_673));
XOR2_X1 i_379 (.Z (n_673), .A (n_659), .B (n_672));
XNOR2_X1 i_378 (.ZN (n_672), .A (n_666), .B (n_671));
XOR2_X1 i_377 (.Z (n_659), .A (n_637), .B (n_658));
XOR2_X1 i_376 (.Z (n_658), .A (n_653), .B (n_657));
XNOR2_X1 i_375 (.ZN (n_657), .A (n_655), .B (n_656));
NAND2_X1 i_374 (.ZN (n_656), .A1 (A[3]), .A2 (B[14]));
XNOR2_X1 i_373 (.ZN (n_655), .A (n_599), .B (n_654));
NAND2_X1 i_372 (.ZN (n_654), .A1 (A[4]), .A2 (B[13]));
XOR2_X1 i_371 (.Z (n_653), .A (n_644), .B (n_652));
XNOR2_X1 i_370 (.ZN (n_652), .A (n_650), .B (n_651));
NAND2_X1 i_369 (.ZN (n_651), .A1 (B[8]), .A2 (A[9]));
OAI21_X1 i_368 (.ZN (n_650), .A (n_649), .B1 (n_646), .B2 (n_648));
NAND2_X1 i_367 (.ZN (n_649), .A1 (n_646), .A2 (n_648));
NOR2_X1 i_366 (.ZN (n_648), .A1 (n_169), .A2 (n_1235));
NOR2_X1 i_365 (.ZN (n_646), .A1 (n_1955), .A2 (n_1339));
XNOR2_X1 i_364 (.ZN (n_644), .A (n_642), .B (n_643));
NAND2_X1 i_363 (.ZN (n_643), .A1 (A[6]), .A2 (B[11]));
NAND2_X1 i_362 (.ZN (n_642), .A1 (n_639), .A2 (n_641));
OAI22_X1 i_361 (.ZN (n_641), .A1 (n_556), .A2 (n_2243), .B1 (n_458), .B2 (n_426));
OR3_X1 i_360 (.ZN (n_639), .A1 (n_638), .A2 (n_556), .A3 (n_426));
NAND2_X1 i_359 (.ZN (n_638), .A1 (B[10]), .A2 (A[8]));
AOI22_X1 i_358 (.ZN (n_637), .A1 (n_595), .A2 (n_596), .B1 (n_636), .B2 (n_594));
INV_X1 i_357 (.ZN (n_636), .A (n_588));
AOI22_X1 i_356 (.ZN (n_635), .A1 (n_618), .A2 (n_619), .B1 (n_597), .B2 (n_617));
OAI21_X1 i_355 (.ZN (n_634), .A (n_633), .B1 (n_628), .B2 (n_632));
NAND2_X1 i_354 (.ZN (n_633), .A1 (n_628), .A2 (n_632));
OAI21_X1 i_353 (.ZN (n_632), .A (n_621), .B1 (n_553), .B2 (n_586));
OAI21_X1 i_352 (.ZN (n_631), .A (n_623), .B1 (n_630), .B2 (n_629));
INV_X1 i_351 (.ZN (n_630), .A (n_624));
XNOR2_X1 i_350 (.ZN (Out[16]), .A (n_625), .B (n_629));
AOI21_X1 i_349 (.ZN (n_629), .A (n_628), .B1 (n_484), .B2 (n_627));
NOR2_X1 i_348 (.ZN (n_628), .A1 (n_484), .A2 (n_627));
INV_X1 i_347 (.ZN (n_627), .A (n_626));
AOI22_X1 i_346 (.ZN (n_626), .A1 (n_510), .A2 (n_547), .B1 (n_486), .B2 (n_509));
NAND2_X1 i_345 (.ZN (n_625), .A1 (n_623), .A2 (n_624));
OR2_X1 i_344 (.ZN (n_624), .A1 (n_551), .A2 (n_622));
NAND2_X1 i_343 (.ZN (n_623), .A1 (n_551), .A2 (n_622));
OAI21_X1 i_342 (.ZN (n_622), .A (n_621), .B1 (n_587), .B2 (n_620));
NAND2_X1 i_341 (.ZN (n_621), .A1 (n_587), .A2 (n_620));
XOR2_X1 i_340 (.Z (n_620), .A (n_618), .B (n_619));
AOI22_X1 i_339 (.ZN (n_619), .A1 (n_507), .A2 (n_508), .B1 (n_505), .B2 (n_506));
XOR2_X1 i_338 (.Z (n_618), .A (n_597), .B (n_617));
XOR2_X1 i_337 (.Z (n_617), .A (n_781), .B (n_782));
XOR2_X1 i_336 (.Z (n_597), .A (n_595), .B (n_596));
AOI22_X1 i_335 (.ZN (n_596), .A1 (n_519), .A2 (n_525), .B1 (n_514), .B2 (n_518));
XNOR2_X1 i_334 (.ZN (n_595), .A (n_588), .B (n_594));
XOR2_X1 i_333 (.Z (n_594), .A (n_576), .B (n_581));
AOI22_X1 i_332 (.ZN (n_588), .A1 (n_500), .A2 (n_504), .B1 (n_493), .B2 (n_499));
XOR2_X1 i_331 (.Z (n_587), .A (n_553), .B (n_586));
XOR2_X1 i_330 (.Z (n_586), .A (n_554), .B (n_585));
XOR2_X1 i_329 (.Z (n_585), .A (n_563), .B (n_584));
XNOR2_X1 i_328 (.ZN (n_584), .A (n_772), .B (n_773));
XNOR2_X1 i_327 (.ZN (n_563), .A (n_495), .B (n_461));
AOI22_X1 i_326 (.ZN (n_554), .A1 (n_539), .A2 (n_545), .B1 (n_529), .B2 (n_538));
AOI22_X1 i_325 (.ZN (n_553), .A1 (n_527), .A2 (n_546), .B1 (n_552), .B2 (n_526));
INV_X1 i_324 (.ZN (n_552), .A (n_512));
INV_X1 i_323 (.ZN (n_551), .A (n_550));
OAI22_X1 i_322 (.ZN (n_550), .A1 (n_479), .A2 (n_549), .B1 (n_485), .B2 (n_548));
XOR2_X1 i_321 (.Z (Out[15]), .A (n_479), .B (n_549));
XNOR2_X1 i_320 (.ZN (n_549), .A (n_485), .B (n_548));
XOR2_X1 i_319 (.Z (n_548), .A (n_510), .B (n_547));
XNOR2_X1 i_318 (.ZN (n_547), .A (n_527), .B (n_546));
XOR2_X1 i_317 (.Z (n_546), .A (n_539), .B (n_545));
XOR2_X1 i_316 (.Z (n_545), .A (n_470), .B (n_462));
XOR2_X1 i_315 (.Z (n_539), .A (n_529), .B (n_538));
XOR2_X1 i_314 (.Z (n_538), .A (n_524), .B (n_516));
AOI22_X1 i_313 (.ZN (n_529), .A1 (n_246), .A2 (n_267), .B1 (n_528), .B2 (n_245));
INV_X1 i_312 (.ZN (n_528), .A (n_222));
XNOR2_X1 i_311 (.ZN (n_527), .A (n_512), .B (n_526));
XNOR2_X1 i_310 (.ZN (n_526), .A (n_519), .B (n_525));
XNOR2_X1 i_309 (.ZN (n_525), .A (n_565), .B (n_566));
XOR2_X1 i_308 (.Z (n_519), .A (n_514), .B (n_518));
XNOR2_X1 i_307 (.ZN (n_518), .A (n_614), .B (n_615));
AOI22_X1 i_306 (.ZN (n_514), .A1 (n_433), .A2 (n_435), .B1 (n_513), .B2 (n_432));
INV_X1 i_305 (.ZN (n_513), .A (n_431));
AOI22_X1 i_304 (.ZN (n_512), .A1 (n_273), .A2 (n_268), .B1 (n_511), .B2 (n_274));
INV_X1 i_303 (.ZN (n_511), .A (n_304));
XOR2_X1 i_302 (.Z (n_510), .A (n_486), .B (n_509));
XOR2_X1 i_301 (.Z (n_509), .A (n_507), .B (n_508));
AOI22_X1 i_300 (.ZN (n_508), .A1 (n_436), .A2 (n_449), .B1 (n_448), .B2 (n_443));
XOR2_X1 i_299 (.Z (n_507), .A (n_505), .B (n_506));
OAI21_X1 i_298 (.ZN (n_506), .A (n_472), .B1 (n_463), .B2 (n_456));
XNOR2_X1 i_297 (.ZN (n_505), .A (n_500), .B (n_504));
XOR2_X1 i_296 (.Z (n_504), .A (n_502), .B (n_503));
NAND2_X1 i_295 (.ZN (n_503), .A1 (A[0]), .A2 (B[15]));
XOR2_X1 i_294 (.Z (n_500), .A (n_493), .B (n_499));
XOR2_X1 i_293 (.Z (n_499), .A (n_497), .B (n_569));
NAND2_X1 i_292 (.ZN (n_497), .A1 (n_571), .A2 (n_568));
XOR2_X1 i_291 (.Z (n_493), .A (n_491), .B (n_579));
NAND2_X1 i_290 (.ZN (n_491), .A1 (n_580), .A2 (n_490));
INV_X1 i_289 (.ZN (n_490), .A (n_578));
OAI21_X1 i_288 (.ZN (n_486), .A (n_451), .B1 (n_452), .B2 (n_473));
OAI21_X1 i_287 (.ZN (n_485), .A (n_484), .B1 (n_480), .B2 (n_483));
NAND2_X1 i_286 (.ZN (n_484), .A1 (n_480), .A2 (n_483));
INV_X1 i_285 (.ZN (n_483), .A (n_482));
AOI22_X1 i_284 (.ZN (n_482), .A1 (n_474), .A2 (n_429), .B1 (n_481), .B2 (n_428));
INV_X1 i_283 (.ZN (n_481), .A (n_415));
INV_X1 i_282 (.ZN (n_480), .A (n_413));
AOI22_X1 i_281 (.ZN (n_479), .A1 (n_477), .A2 (n_476), .B1 (n_478), .B2 (n_475));
INV_X1 i_280 (.ZN (n_478), .A (n_414));
XOR2_X1 i_279 (.Z (Out[14]), .A (n_476), .B (n_477));
OAI22_X1 i_278 (.ZN (n_477), .A1 (n_409), .A2 (n_407), .B1 (n_366), .B2 (n_406));
XNOR2_X1 i_277 (.ZN (n_476), .A (n_414), .B (n_475));
XOR2_X1 i_276 (.Z (n_475), .A (n_429), .B (n_474));
XNOR2_X1 i_275 (.ZN (n_474), .A (n_452), .B (n_473));
OAI21_X1 i_274 (.ZN (n_473), .A (n_472), .B1 (n_464), .B2 (n_471));
NAND2_X1 i_273 (.ZN (n_472), .A1 (n_464), .A2 (n_471));
XNOR2_X1 i_272 (.ZN (n_471), .A (n_541), .B (n_540));
XOR2_X1 i_271 (.Z (n_464), .A (n_456), .B (n_463));
XOR2_X1 i_270 (.Z (n_463), .A (n_466), .B (n_465));
XOR2_X1 i_269 (.Z (n_456), .A (n_492), .B (n_489));
OAI21_X1 i_268 (.ZN (n_452), .A (n_451), .B1 (n_430), .B2 (n_450));
NAND2_X1 i_267 (.ZN (n_451), .A1 (n_430), .A2 (n_450));
XNOR2_X1 i_266 (.ZN (n_450), .A (n_436), .B (n_449));
XOR2_X1 i_265 (.Z (n_449), .A (n_443), .B (n_448));
XNOR2_X1 i_264 (.ZN (n_448), .A (n_447), .B (n_287));
NOR2_X1 i_263 (.ZN (n_447), .A1 (n_534), .A2 (n_537));
XOR2_X1 i_262 (.Z (n_443), .A (n_440), .B (n_517));
NOR2_X1 i_261 (.ZN (n_440), .A1 (n_520), .A2 (n_523));
XOR2_X1 i_260 (.Z (n_436), .A (n_433), .B (n_435));
AOI21_X1 i_259 (.ZN (n_435), .A (n_285), .B1 (n_434), .B2 (n_284));
INV_X1 i_258 (.ZN (n_434), .A (n_286));
XNOR2_X1 i_257 (.ZN (n_433), .A (n_431), .B (n_432));
AOI21_X1 i_256 (.ZN (n_432), .A (n_281), .B1 (n_283), .B2 (n_270));
AOI21_X1 i_255 (.ZN (n_431), .A (n_309), .B1 (n_307), .B2 (n_306));
AOI22_X1 i_254 (.ZN (n_430), .A1 (n_361), .A2 (n_362), .B1 (n_353), .B2 (n_360));
XNOR2_X1 i_253 (.ZN (n_429), .A (n_415), .B (n_428));
XOR2_X1 i_252 (.Z (n_428), .A (n_273), .B (n_268));
AOI22_X1 i_251 (.ZN (n_415), .A1 (n_403), .A2 (n_402), .B1 (n_383), .B2 (n_401));
OAI21_X1 i_250 (.ZN (n_414), .A (n_413), .B1 (n_411), .B2 (n_412));
NAND2_X1 i_249 (.ZN (n_413), .A1 (n_411), .A2 (n_412));
INV_X1 i_248 (.ZN (n_412), .A (n_405));
AOI22_X1 i_247 (.ZN (n_411), .A1 (n_365), .A2 (n_364), .B1 (n_410), .B2 (n_363));
INV_X1 i_246 (.ZN (n_410), .A (n_352));
XOR2_X1 i_245 (.Z (Out[13]), .A (n_407), .B (n_409));
AOI22_X1 i_244 (.ZN (n_409), .A1 (n_351), .A2 (n_348), .B1 (n_408), .B2 (n_344));
INV_X1 i_243 (.ZN (n_408), .A (n_347));
XNOR2_X1 i_242 (.ZN (n_407), .A (n_366), .B (n_406));
OAI21_X1 i_241 (.ZN (n_406), .A (n_405), .B1 (n_367), .B2 (n_404));
NAND2_X1 i_240 (.ZN (n_405), .A1 (n_367), .A2 (n_404));
XOR2_X1 i_239 (.Z (n_404), .A (n_402), .B (n_403));
AOI22_X1 i_238 (.ZN (n_403), .A1 (n_303), .A2 (n_316), .B1 (n_310), .B2 (n_315));
XOR2_X1 i_237 (.Z (n_402), .A (n_383), .B (n_401));
XNOR2_X1 i_236 (.ZN (n_401), .A (n_276), .B (n_275));
XOR2_X1 i_235 (.Z (n_383), .A (n_312), .B (n_305));
INV_X1 i_234 (.ZN (n_367), .A (n_346));
XOR2_X1 i_233 (.Z (n_366), .A (n_364), .B (n_365));
AOI22_X1 i_232 (.ZN (n_365), .A1 (n_318), .A2 (n_343), .B1 (n_296), .B2 (n_317));
XNOR2_X1 i_231 (.ZN (n_364), .A (n_352), .B (n_363));
XNOR2_X1 i_230 (.ZN (n_363), .A (n_361), .B (n_362));
AOI22_X1 i_229 (.ZN (n_362), .A1 (n_337), .A2 (n_341), .B1 (n_329), .B2 (n_336));
XOR2_X1 i_228 (.Z (n_361), .A (n_353), .B (n_360));
XOR2_X1 i_227 (.Z (n_360), .A (n_189), .B (n_212));
OAI22_X1 i_226 (.ZN (n_353), .A1 (n_298), .A2 (n_302), .B1 (n_300), .B2 (n_301));
AOI22_X1 i_225 (.ZN (n_352), .A1 (n_322), .A2 (n_342), .B1 (n_427), .B2 (n_354));
XOR2_X1 i_224 (.Z (Out[12]), .A (n_348), .B (n_351));
AOI22_X1 i_223 (.ZN (n_351), .A1 (n_349), .A2 (n_294), .B1 (n_350), .B2 (n_290));
INV_X1 i_222 (.ZN (n_350), .A (n_293));
INV_X1 i_221 (.ZN (n_349), .A (n_295));
XNOR2_X1 i_220 (.ZN (n_348), .A (n_344), .B (n_347));
OAI21_X1 i_219 (.ZN (n_347), .A (n_346), .B1 (n_292), .B2 (n_345));
NAND2_X1 i_218 (.ZN (n_346), .A1 (n_345), .A2 (n_292));
OAI22_X1 i_217 (.ZN (n_345), .A1 (n_255), .A2 (n_289), .B1 (n_271), .B2 (n_288));
XOR2_X1 i_216 (.Z (n_344), .A (n_318), .B (n_343));
XNOR2_X1 i_215 (.ZN (n_343), .A (n_322), .B (n_342));
XOR2_X1 i_214 (.Z (n_342), .A (n_337), .B (n_341));
XNOR2_X1 i_213 (.ZN (n_341), .A (n_177), .B (n_178));
XOR2_X1 i_212 (.Z (n_337), .A (n_329), .B (n_336));
OAI21_X1 i_211 (.ZN (n_336), .A (n_174), .B1 (n_168), .B2 (n_171));
XNOR2_X1 i_210 (.ZN (n_329), .A (n_262), .B (n_263));
XOR2_X1 i_209 (.Z (n_322), .A (n_427), .B (n_354));
XOR2_X1 i_208 (.Z (n_318), .A (n_296), .B (n_317));
XNOR2_X1 i_207 (.ZN (n_317), .A (n_303), .B (n_316));
XOR2_X1 i_206 (.Z (n_316), .A (n_310), .B (n_315));
XOR2_X1 i_205 (.Z (n_315), .A (n_207), .B (n_208));
XNOR2_X1 i_204 (.ZN (n_310), .A (n_321), .B (n_269));
XNOR2_X1 i_203 (.ZN (n_303), .A (n_298), .B (n_302));
XNOR2_X1 i_202 (.ZN (n_302), .A (n_300), .B (n_301));
AOI21_X1 i_201 (.ZN (n_301), .A (n_369), .B1 (n_359), .B2 (n_358));
AOI21_X1 i_200 (.ZN (n_300), .A (n_373), .B1 (n_371), .B2 (n_299));
INV_X1 i_199 (.ZN (n_299), .A (n_198));
AOI22_X1 i_198 (.ZN (n_298), .A1 (n_249), .A2 (n_250), .B1 (n_247), .B2 (n_297));
INV_X1 i_197 (.ZN (n_297), .A (n_248));
AOI22_X1 i_196 (.ZN (n_296), .A1 (n_252), .A2 (n_254), .B1 (n_244), .B2 (n_251));
XOR2_X1 i_195 (.Z (Out[11]), .A (n_294), .B (n_295));
AOI22_X1 i_194 (.ZN (n_295), .A1 (n_243), .A2 (n_242), .B1 (n_235), .B2 (n_241));
XNOR2_X1 i_193 (.ZN (n_294), .A (n_290), .B (n_293));
AOI21_X1 i_192 (.ZN (n_293), .A (n_292), .B1 (n_240), .B2 (n_291));
NOR2_X1 i_191 (.ZN (n_292), .A1 (n_291), .A2 (n_240));
OAI21_X1 i_190 (.ZN (n_291), .A (n_220), .B1 (n_221), .B2 (n_234));
XNOR2_X1 i_189 (.ZN (n_290), .A (n_255), .B (n_289));
XNOR2_X1 i_188 (.ZN (n_289), .A (n_271), .B (n_288));
XNOR2_X1 i_187 (.ZN (n_288), .A (n_375), .B (n_355));
XNOR2_X1 i_186 (.ZN (n_271), .A (n_439), .B (n_437));
XOR2_X1 i_185 (.Z (n_255), .A (n_252), .B (n_254));
AOI22_X1 i_184 (.ZN (n_254), .A1 (n_232), .A2 (n_253), .B1 (n_231), .B2 (n_225));
INV_X1 i_183 (.ZN (n_253), .A (n_233));
XOR2_X1 i_182 (.Z (n_252), .A (n_244), .B (n_251));
XNOR2_X1 i_181 (.ZN (n_251), .A (n_249), .B (n_250));
OAI22_X1 i_180 (.ZN (n_250), .A1 (n_224), .A2 (n_385), .B1 (n_374), .B2 (n_223));
XNOR2_X1 i_179 (.ZN (n_249), .A (n_247), .B (n_248));
AOI21_X1 i_178 (.ZN (n_248), .A (n_199), .B1 (n_201), .B2 (n_202));
OAI33_X1 i_177 (.ZN (n_247), .A1 (n_214), .A2 (n_99), .A3 (n_1955), .B1 (n_389), .B2 (n_423), .B3 (n_169));
AOI22_X1 i_176 (.ZN (n_244), .A1 (n_211), .A2 (n_216), .B1 (n_210), .B2 (n_203));
XNOR2_X1 i_175 (.ZN (Out[10]), .A (n_242), .B (n_243));
OAI21_X1 i_174 (.ZN (n_243), .A (n_196), .B1 (n_160), .B2 (n_197));
XOR2_X1 i_173 (.Z (n_242), .A (n_235), .B (n_241));
OAI21_X1 i_172 (.ZN (n_241), .A (n_240), .B1 (n_236), .B2 (n_239));
NAND2_X1 i_171 (.ZN (n_240), .A1 (n_236), .A2 (n_239));
AOI21_X1 i_170 (.ZN (n_239), .A (n_237), .B1 (n_180), .B2 (n_238));
INV_X1 i_169 (.ZN (n_238), .A (n_194));
INV_X1 i_168 (.ZN (n_237), .A (n_193));
INV_X1 i_167 (.ZN (n_236), .A (n_162));
XOR2_X1 i_166 (.Z (n_235), .A (n_221), .B (n_234));
XNOR2_X1 i_165 (.ZN (n_234), .A (n_232), .B (n_233));
AOI22_X1 i_164 (.ZN (n_233), .A1 (n_186), .A2 (n_190), .B1 (n_184), .B2 (n_185));
XOR2_X1 i_163 (.Z (n_232), .A (n_225), .B (n_231));
XOR2_X1 i_162 (.Z (n_231), .A (n_376), .B (n_390));
XOR2_X1 i_161 (.Z (n_225), .A (n_224), .B (n_385));
XNOR2_X1 i_160 (.ZN (n_224), .A (n_374), .B (n_223));
NAND2_X1 i_159 (.ZN (n_223), .A1 (A[0]), .A2 (B[10]));
OAI21_X1 i_158 (.ZN (n_221), .A (n_220), .B1 (n_217), .B2 (n_219));
NAND2_X1 i_157 (.ZN (n_220), .A1 (n_217), .A2 (n_219));
OAI22_X1 i_156 (.ZN (n_219), .A1 (n_173), .A2 (n_179), .B1 (n_218), .B2 (n_172));
INV_X1 i_155 (.ZN (n_218), .A (n_165));
XNOR2_X1 i_154 (.ZN (n_217), .A (n_211), .B (n_216));
XOR2_X1 i_153 (.Z (n_216), .A (n_214), .B (n_215));
NAND2_X1 i_152 (.ZN (n_215), .A1 (A[3]), .A2 (B[7]));
XNOR2_X1 i_151 (.ZN (n_214), .A (n_370), .B (n_213));
NAND2_X1 i_150 (.ZN (n_213), .A1 (B[5]), .A2 (A[5]));
XOR2_X1 i_149 (.Z (n_211), .A (n_203), .B (n_210));
XOR2_X1 i_148 (.Z (n_210), .A (n_446), .B (n_445));
XOR2_X1 i_147 (.Z (n_203), .A (n_201), .B (n_202));
NOR2_X1 i_146 (.ZN (n_202), .A1 (n_340), .A2 (n_170));
NOR2_X1 i_145 (.ZN (n_201), .A1 (n_199), .A2 (n_200));
AOI22_X1 i_144 (.ZN (n_200), .A1 (B[3]), .A2 (A[7]), .B1 (B[2]), .B2 (A[8]));
NOR2_X1 i_143 (.ZN (n_199), .A1 (n_455), .A2 (n_331));
XNOR2_X1 i_142 (.ZN (Out[9]), .A (n_160), .B (n_197));
OAI21_X1 i_141 (.ZN (n_197), .A (n_196), .B1 (n_163), .B2 (n_195));
NAND2_X1 i_140 (.ZN (n_196), .A1 (n_163), .A2 (n_195));
XNOR2_X1 i_139 (.ZN (n_195), .A (n_180), .B (n_194));
OAI21_X1 i_138 (.ZN (n_194), .A (n_193), .B1 (n_191), .B2 (n_192));
NAND2_X1 i_137 (.ZN (n_193), .A1 (n_191), .A2 (n_192));
OAI22_X1 i_136 (.ZN (n_192), .A1 (n_145), .A2 (n_152), .B1 (n_144), .B2 (n_138));
XNOR2_X1 i_135 (.ZN (n_191), .A (n_186), .B (n_190));
XOR2_X1 i_134 (.Z (n_190), .A (n_388), .B (n_387));
XOR2_X1 i_133 (.Z (n_186), .A (n_184), .B (n_185));
OAI22_X1 i_132 (.ZN (n_185), .A1 (n_136), .A2 (n_137), .B1 (n_386), .B2 (n_135));
XOR2_X1 i_131 (.Z (n_184), .A (n_454), .B (n_183));
NAND2_X1 i_130 (.ZN (n_183), .A1 (B[3]), .A2 (A[6]));
XOR2_X1 i_129 (.Z (n_180), .A (n_173), .B (n_179));
XOR2_X1 i_128 (.Z (n_179), .A (n_397), .B (n_391));
XOR2_X1 i_127 (.Z (n_173), .A (n_165), .B (n_172));
XOR2_X1 i_126 (.Z (n_172), .A (n_381), .B (n_380));
AOI22_X1 i_125 (.ZN (n_165), .A1 (n_128), .A2 (n_129), .B1 (n_125), .B2 (n_164));
INV_X1 i_124 (.ZN (n_164), .A (n_127));
OAI21_X1 i_123 (.ZN (n_163), .A (n_162), .B1 (n_161), .B2 (n_154));
NAND2_X1 i_122 (.ZN (n_162), .A1 (n_161), .A2 (n_154));
AOI22_X1 i_121 (.ZN (n_161), .A1 (n_131), .A2 (n_105), .B1 (n_124), .B2 (n_130));
AOI21_X1 i_120 (.ZN (n_160), .A (n_158), .B1 (n_123), .B2 (n_156));
XNOR2_X1 i_119 (.ZN (Out[8]), .A (n_123), .B (n_159));
NOR2_X1 i_118 (.ZN (n_159), .A1 (n_157), .A2 (n_158));
NOR2_X1 i_117 (.ZN (n_158), .A1 (n_132), .A2 (n_155));
INV_X1 i_116 (.ZN (n_157), .A (n_156));
NAND2_X1 i_115 (.ZN (n_156), .A1 (n_132), .A2 (n_155));
AOI21_X1 i_114 (.ZN (n_155), .A (n_154), .B1 (n_134), .B2 (n_153));
NOR2_X1 i_113 (.ZN (n_154), .A1 (n_134), .A2 (n_153));
XOR2_X1 i_112 (.Z (n_153), .A (n_145), .B (n_152));
XOR2_X1 i_111 (.Z (n_152), .A (n_393), .B (n_392));
XNOR2_X1 i_110 (.ZN (n_145), .A (n_138), .B (n_144));
XOR2_X1 i_109 (.Z (n_144), .A (n_417), .B (n_416));
XOR2_X1 i_108 (.Z (n_138), .A (n_136), .B (n_137));
NAND2_X1 i_107 (.ZN (n_137), .A1 (A[0]), .A2 (B[8]));
XNOR2_X1 i_106 (.ZN (n_136), .A (n_386), .B (n_135));
NAND2_X1 i_105 (.ZN (n_135), .A1 (A[2]), .A2 (B[6]));
AOI22_X1 i_104 (.ZN (n_134), .A1 (n_133), .A2 (n_118), .B1 (n_111), .B2 (n_117));
INV_X1 i_103 (.ZN (n_133), .A (n_88));
XNOR2_X1 i_102 (.ZN (n_132), .A (n_131), .B (n_105));
XOR2_X1 i_101 (.Z (n_131), .A (n_124), .B (n_130));
XNOR2_X1 i_100 (.ZN (n_130), .A (n_128), .B (n_129));
OAI22_X1 i_99 (.ZN (n_129), .A1 (n_98), .A2 (n_101), .B1 (n_421), .B2 (n_100));
XNOR2_X1 i_98 (.ZN (n_128), .A (n_125), .B (n_127));
AOI21_X1 i_97 (.ZN (n_127), .A (n_108), .B1 (n_110), .B2 (n_126));
INV_X1 i_96 (.ZN (n_126), .A (n_71));
OAI21_X1 i_95 (.ZN (n_125), .A (n_114), .B1 (n_116), .B2 (n_112));
AOI22_X1 i_94 (.ZN (n_124), .A1 (n_97), .A2 (n_102), .B1 (n_93), .B2 (n_96));
AOI22_X1 i_93 (.ZN (n_123), .A1 (n_120), .A2 (n_121), .B1 (n_122), .B2 (n_119));
INV_X1 i_92 (.ZN (n_122), .A (n_106));
XOR2_X1 i_91 (.Z (Out[7]), .A (n_120), .B (n_121));
AOI22_X1 i_90 (.ZN (n_121), .A1 (n_90), .A2 (n_91), .B1 (n_85), .B2 (n_89));
XNOR2_X1 i_89 (.ZN (n_120), .A (n_106), .B (n_119));
XNOR2_X1 i_88 (.ZN (n_119), .A (n_88), .B (n_118));
XOR2_X1 i_87 (.Z (n_118), .A (n_111), .B (n_117));
XOR2_X1 i_86 (.Z (n_117), .A (n_112), .B (n_116));
NAND2_X1 i_85 (.ZN (n_116), .A1 (n_114), .A2 (n_115));
OAI21_X1 i_84 (.ZN (n_115), .A (n_77), .B1 (n_424), .B2 (n_422));
OR3_X1 i_83 (.ZN (n_114), .A1 (n_77), .A2 (n_424), .A3 (n_422));
NAND2_X1 i_82 (.ZN (n_112), .A1 (B[4]), .A2 (A[3]));
XNOR2_X1 i_81 (.ZN (n_111), .A (n_110), .B (n_71));
NOR2_X1 i_80 (.ZN (n_110), .A1 (n_108), .A2 (n_109));
AOI22_X1 i_79 (.ZN (n_109), .A1 (A[1]), .A2 (B[6]), .B1 (A[0]), .B2 (B[7]));
NOR2_X1 i_78 (.ZN (n_108), .A1 (n_75), .A2 (n_386));
OAI21_X1 i_77 (.ZN (n_106), .A (n_105), .B1 (n_103), .B2 (n_104));
NAND2_X1 i_76 (.ZN (n_105), .A1 (n_103), .A2 (n_104));
OAI21_X1 i_75 (.ZN (n_104), .A (n_83), .B1 (n_70), .B2 (n_84));
XOR2_X1 i_74 (.Z (n_103), .A (n_97), .B (n_102));
XOR2_X1 i_73 (.Z (n_102), .A (n_98), .B (n_101));
XNOR2_X1 i_72 (.ZN (n_101), .A (n_421), .B (n_100));
NAND2_X1 i_71 (.ZN (n_100), .A1 (B[1]), .A2 (A[6]));
AOI21_X1 i_70 (.ZN (n_98), .A (n_78), .B1 (n_80), .B2 (n_81));
OAI22_X1 i_69 (.ZN (n_97), .A1 (n_93), .A2 (n_95), .B1 (n_92), .B2 (n_96));
INV_X1 i_68 (.ZN (n_96), .A (n_95));
AOI21_X1 i_67 (.ZN (n_95), .A (n_72), .B1 (n_74), .B2 (n_94));
INV_X1 i_66 (.ZN (n_94), .A (n_75));
INV_X1 i_65 (.ZN (n_93), .A (n_92));
AOI22_X1 i_64 (.ZN (n_92), .A1 (n_68), .A2 (n_69), .B1 (n_67), .B2 (n_65));
XNOR2_X1 i_63 (.ZN (Out[6]), .A (n_90), .B (n_91));
OAI22_X1 i_62 (.ZN (n_91), .A1 (n_62), .A2 (n_63), .B1 (n_56), .B2 (n_61));
XOR2_X1 i_61 (.Z (n_90), .A (n_85), .B (n_89));
NAND2_X1 i_60 (.ZN (n_89), .A1 (n_87), .A2 (n_88));
OR3_X1 i_59 (.ZN (n_88), .A1 (n_86), .A2 (n_46), .A3 (n_60));
OAI21_X1 i_58 (.ZN (n_87), .A (n_86), .B1 (n_46), .B2 (n_60));
AOI22_X1 i_57 (.ZN (n_86), .A1 (n_51), .A2 (n_55), .B1 (n_50), .B2 (n_42));
XNOR2_X1 i_56 (.ZN (n_85), .A (n_70), .B (n_84));
OAI21_X1 i_55 (.ZN (n_84), .A (n_83), .B1 (n_76), .B2 (n_82));
NAND2_X1 i_54 (.ZN (n_83), .A1 (n_76), .A2 (n_82));
XOR2_X1 i_53 (.Z (n_82), .A (n_80), .B (n_81));
NOR2_X1 i_52 (.ZN (n_81), .A1 (n_424), .A2 (n_99));
NOR2_X1 i_51 (.ZN (n_80), .A1 (n_78), .A2 (n_79));
AOI22_X1 i_50 (.ZN (n_79), .A1 (B[2]), .A2 (A[4]), .B1 (B[1]), .B2 (A[5]));
NOR2_X1 i_49 (.ZN (n_78), .A1 (n_39), .A2 (n_77));
NAND2_X1 i_48 (.ZN (n_77), .A1 (B[2]), .A2 (A[5]));
XNOR2_X1 i_47 (.ZN (n_76), .A (n_74), .B (n_75));
NAND2_X1 i_46 (.ZN (n_75), .A1 (A[0]), .A2 (B[6]));
NOR2_X1 i_45 (.ZN (n_74), .A1 (n_72), .A2 (n_73));
AOI22_X1 i_44 (.ZN (n_73), .A1 (A[2]), .A2 (B[4]), .B1 (A[1]), .B2 (B[5]));
NOR2_X1 i_43 (.ZN (n_72), .A1 (n_57), .A2 (n_71));
NAND2_X1 i_42 (.ZN (n_71), .A1 (A[2]), .A2 (B[5]));
XNOR2_X1 i_41 (.ZN (n_70), .A (n_68), .B (n_69));
OAI22_X1 i_40 (.ZN (n_69), .A1 (n_58), .A2 (n_59), .B1 (n_30), .B2 (n_57));
XOR2_X1 i_39 (.Z (n_68), .A (n_65), .B (n_67));
OAI33_X1 i_38 (.ZN (n_67), .A1 (n_53), .A2 (n_29), .A3 (n_99), .B1 (n_39), .B2 (n_28), .B3 (n_423));
NOR2_X1 i_37 (.ZN (n_65), .A1 (n_28), .A2 (n_170));
XNOR2_X1 i_36 (.ZN (Out[5]), .A (n_62), .B (n_63));
AOI22_X1 i_35 (.ZN (n_63), .A1 (n_48), .A2 (n_49), .B1 (n_47), .B2 (n_37));
XNOR2_X1 i_34 (.ZN (n_62), .A (n_56), .B (n_61));
XOR2_X1 i_33 (.Z (n_61), .A (n_60), .B (n_46));
XNOR2_X1 i_32 (.ZN (n_60), .A (n_58), .B (n_59));
NAND2_X1 i_31 (.ZN (n_59), .A1 (A[0]), .A2 (B[5]));
XNOR2_X1 i_30 (.ZN (n_58), .A (n_30), .B (n_57));
NAND2_X1 i_29 (.ZN (n_57), .A1 (A[1]), .A2 (B[4]));
XOR2_X1 i_28 (.Z (n_56), .A (n_51), .B (n_55));
XOR2_X1 i_27 (.Z (n_55), .A (n_53), .B (n_54));
NAND2_X1 i_26 (.ZN (n_54), .A1 (B[2]), .A2 (A[3]));
XNOR2_X1 i_25 (.ZN (n_53), .A (n_39), .B (n_52));
NAND2_X1 i_24 (.ZN (n_52), .A1 (B[0]), .A2 (A[5]));
XNOR2_X1 i_23 (.ZN (n_51), .A (n_50), .B (n_41));
OAI21_X1 i_22 (.ZN (n_50), .A (n_32), .B1 (n_35), .B2 (n_36));
XNOR2_X1 i_21 (.ZN (Out[4]), .A (n_48), .B (n_49));
OAI21_X1 i_20 (.ZN (n_49), .A (n_143), .B1 (n_141), .B2 (n_149));
XOR2_X1 i_19 (.Z (n_48), .A (n_37), .B (n_47));
OAI21_X1 i_18 (.ZN (n_47), .A (n_46), .B1 (n_44), .B2 (n_45));
NAND2_X1 i_17 (.ZN (n_46), .A1 (n_44), .A2 (n_45));
AOI21_X1 i_16 (.ZN (n_45), .A (n_66), .B1 (n_150), .B2 (n_64));
OAI21_X1 i_15 (.ZN (n_44), .A (n_38), .B1 (n_42), .B2 (n_43));
AOI22_X1 i_14 (.ZN (n_43), .A1 (B[0]), .A2 (A[4]), .B1 (B[1]), .B2 (A[3]));
INV_X1 i_13 (.ZN (n_42), .A (n_41));
OAI21_X1 i_12 (.ZN (n_41), .A (n_107), .B1 (n_25), .B2 (n_40));
INV_X1 i_11 (.ZN (n_40), .A (n_39));
NAND2_X1 i_10 (.ZN (n_39), .A1 (B[1]), .A2 (A[4]));
NAND3_X1 i_9 (.ZN (n_38), .A1 (n_25), .A2 (A[4]), .A3 (n_107));
XNOR2_X1 i_8 (.ZN (n_37), .A (n_35), .B (n_36));
NAND2_X1 i_7 (.ZN (n_36), .A1 (A[0]), .A2 (B[4]));
NAND2_X1 i_6 (.ZN (n_35), .A1 (n_32), .A2 (n_34));
OAI22_X1 i_5 (.ZN (n_34), .A1 (n_1534), .A2 (n_424), .B1 (n_29), .B2 (n_33));
OR3_X1 i_4 (.ZN (n_32), .A1 (n_30), .A2 (n_1534), .A3 (n_29));
NAND2_X1 i_3 (.ZN (n_30), .A1 (A[2]), .A2 (B[3]));
NOR2_X1 i_2 (.ZN (Out[1]), .A1 (n_19), .A2 (n_3));
AOI22_X1 i_1 (.ZN (n_3), .A1 (A[0]), .A2 (B[1]), .B1 (B[0]), .B2 (A[1]));
INV_X1 i_0 (.ZN (Out[0]), .A (n_20));

endmodule //datapath

module N_Bit_Mult (A, B, Out);

output [47:0] Out;
input [23:0] A;
input [23:0] B;


datapath i_0 (.Out ({Out[47], Out[46], Out[45], Out[44], Out[43], Out[42], Out[41], 
    Out[40], Out[39], Out[38], Out[37], Out[36], Out[35], Out[34], Out[33], Out[32], 
    Out[31], Out[30], Out[29], Out[28], Out[27], Out[26], Out[25], Out[24], Out[23], 
    Out[22], Out[21], Out[20], Out[19], Out[18], Out[17], Out[16], Out[15], Out[14], 
    Out[13], Out[12], Out[11], Out[10], Out[9], Out[8], Out[7], Out[6], Out[5], Out[4], 
    Out[3], Out[2], Out[1], Out[0]}), .A ({A[23], A[22], A[21], A[20], A[19], A[18], 
    A[17], A[16], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], 
    A[5], A[4], A[3], A[2], A[1], A[0]}), .B ({B[23], B[22], B[21], B[20], B[19], 
    B[18], B[17], B[16], B[15], B[14], B[13], B[12], B[11], B[10], B[9], B[8], B[7], 
    B[6], B[5], B[4], B[3], B[2], B[1], B[0]}));

endmodule //N_Bit_Mult

module Reg__0_18 (in, clk, out);

output [31:0] out;
input clk;
input [31:0] in;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk), .D (in[0]));
DFF_X2 \out_reg[1]  (.Q (out[1]), .CK (clk), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk), .D (in[7]));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (clk), .D (in[8]));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (clk), .D (in[9]));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (clk), .D (in[10]));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (clk), .D (in[11]));
DFF_X2 \out_reg[12]  (.Q (out[12]), .CK (clk), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk), .D (in[13]));
DFF_X2 \out_reg[14]  (.Q (out[14]), .CK (clk), .D (in[14]));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (clk), .D (in[15]));
DFF_X2 \out_reg[16]  (.Q (out[16]), .CK (clk), .D (in[16]));
DFF_X2 \out_reg[17]  (.Q (out[17]), .CK (clk), .D (in[17]));
DFF_X2 \out_reg[18]  (.Q (out[18]), .CK (clk), .D (in[18]));
DFF_X2 \out_reg[19]  (.Q (out[19]), .CK (clk), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk), .D (in[20]));
DFF_X2 \out_reg[21]  (.Q (out[21]), .CK (clk), .D (in[21]));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (clk), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk), .D (in[31]));

endmodule //Reg__0_18

module Reg__0_17 (in, clk, out);

output [31:0] out;
input clk;
input [31:0] in;


DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (clk), .D (in[0]));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (clk), .D (in[1]));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (clk), .D (in[2]));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (clk), .D (in[3]));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (clk), .D (in[4]));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (clk), .D (in[5]));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (clk), .D (in[6]));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (clk), .D (in[7]));
DFF_X2 \out_reg[8]  (.Q (out[8]), .CK (clk), .D (in[8]));
DFF_X2 \out_reg[9]  (.Q (out[9]), .CK (clk), .D (in[9]));
DFF_X2 \out_reg[10]  (.Q (out[10]), .CK (clk), .D (in[10]));
DFF_X2 \out_reg[11]  (.Q (out[11]), .CK (clk), .D (in[11]));
DFF_X2 \out_reg[12]  (.Q (out[12]), .CK (clk), .D (in[12]));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (clk), .D (in[13]));
DFF_X2 \out_reg[14]  (.Q (out[14]), .CK (clk), .D (in[14]));
DFF_X2 \out_reg[15]  (.Q (out[15]), .CK (clk), .D (in[15]));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (clk), .D (in[16]));
DFF_X2 \out_reg[17]  (.Q (out[17]), .CK (clk), .D (in[17]));
DFF_X2 \out_reg[18]  (.Q (out[18]), .CK (clk), .D (in[18]));
DFF_X2 \out_reg[19]  (.Q (out[19]), .CK (clk), .D (in[19]));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (clk), .D (in[20]));
DFF_X2 \out_reg[21]  (.Q (out[21]), .CK (clk), .D (in[21]));
DFF_X2 \out_reg[22]  (.Q (out[22]), .CK (clk), .D (in[22]));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (clk), .D (in[23]));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (clk), .D (in[24]));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (clk), .D (in[25]));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (clk), .D (in[26]));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (clk), .D (in[27]));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (clk), .D (in[28]));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (clk), .D (in[29]));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (clk), .D (in[30]));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (clk), .D (in[31]));

endmodule //Reg__0_17

module float_mult (A, B, clk, Exception, Overflow, Underflow, Out);

output Exception;
output [31:0] Out;
output Overflow;
output Underflow;
input [31:0] A;
input [31:0] B;
input clk;
wire \afterB[31] ;
wire \afterB[30] ;
wire \afterB[29] ;
wire \afterB[28] ;
wire \afterB[27] ;
wire \afterB[26] ;
wire \afterB[25] ;
wire \afterB[24] ;
wire \afterB[23] ;
wire \afterB[22] ;
wire \afterB[21] ;
wire \afterB[20] ;
wire \afterB[19] ;
wire \afterB[18] ;
wire \afterB[17] ;
wire \afterB[16] ;
wire \afterB[15] ;
wire \afterB[14] ;
wire \afterB[13] ;
wire \afterB[12] ;
wire \afterB[11] ;
wire \afterB[10] ;
wire \afterB[9] ;
wire \afterB[8] ;
wire \afterB[7] ;
wire \afterB[6] ;
wire \afterB[5] ;
wire \afterB[4] ;
wire \afterB[3] ;
wire \afterB[2] ;
wire \afterB[1] ;
wire \afterB[0] ;
wire \afterA[31] ;
wire \afterA[30] ;
wire \afterA[29] ;
wire \afterA[28] ;
wire \afterA[27] ;
wire \afterA[26] ;
wire \afterA[25] ;
wire \afterA[24] ;
wire \afterA[23] ;
wire \afterA[22] ;
wire \afterA[21] ;
wire \afterA[20] ;
wire \afterA[19] ;
wire \afterA[18] ;
wire \afterA[17] ;
wire \afterA[16] ;
wire \afterA[15] ;
wire \afterA[14] ;
wire \afterA[13] ;
wire \afterA[12] ;
wire \afterA[11] ;
wire \afterA[10] ;
wire \afterA[9] ;
wire \afterA[8] ;
wire \afterA[7] ;
wire \afterA[6] ;
wire \afterA[5] ;
wire \afterA[4] ;
wire \afterA[3] ;
wire \afterA[2] ;
wire \afterA[1] ;
wire \afterA[0] ;
wire \MP[47] ;
wire \MP[46] ;
wire \MP[45] ;
wire \MP[44] ;
wire \MP[43] ;
wire \MP[42] ;
wire \MP[41] ;
wire \MP[40] ;
wire \MP[39] ;
wire \MP[38] ;
wire \MP[37] ;
wire \MP[36] ;
wire \MP[35] ;
wire \MP[34] ;
wire \MP[33] ;
wire \MP[32] ;
wire \MP[31] ;
wire \MP[30] ;
wire \MP[29] ;
wire \MP[28] ;
wire \MP[27] ;
wire \MP[26] ;
wire \MP[25] ;
wire \MP[24] ;
wire \MP[23] ;
wire \MP[22] ;
wire \MP[21] ;
wire \MP[20] ;
wire \MP[19] ;
wire \MP[18] ;
wire \MP[17] ;
wire \MP[16] ;
wire \MP[15] ;
wire \MP[14] ;
wire \MP[13] ;
wire \MP[12] ;
wire \MP[11] ;
wire \MP[10] ;
wire \MP[9] ;
wire \MP[8] ;
wire \MP[7] ;
wire \MP[6] ;
wire \MP[5] ;
wire \MP[4] ;
wire \MP[3] ;
wire \MP[2] ;
wire \MP[1] ;
wire \MP[0] ;
wire \MP_final[22] ;
wire \MP_final[21] ;
wire \MP_final[20] ;
wire \MP_final[19] ;
wire \MP_final[18] ;
wire \MP_final[17] ;
wire \MP_final[16] ;
wire \MP_final[15] ;
wire \MP_final[14] ;
wire \MP_final[13] ;
wire \MP_final[12] ;
wire \MP_final[11] ;
wire \MP_final[10] ;
wire \MP_final[9] ;
wire \MP_final[8] ;
wire \MP_final[7] ;
wire \MP_final[6] ;
wire \MP_final[5] ;
wire \MP_final[4] ;
wire \MP_final[3] ;
wire \MP_final[2] ;
wire \MP_final[1] ;
wire \MP_final[0] ;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_0_0;
wire n_0_23;
wire n_0_0_1;
wire n_0_0_2;
wire n_0_24;
wire n_0_25;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_26;
wire n_0_0_7;
wire n_0_27;
wire n_0_0_8;
wire n_0_28;
wire n_0_29;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_30;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_31;
wire n_0_0_15;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_0_39;
wire n_0_0_41;
wire n_0_0_42;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire n_0_0_71;
wire n_0_0_72;
wire n_0_0_73;
wire n_0_0_74;
wire n_0_0_75;
wire n_0_34;
wire n_0_0_79;
wire n_0_0_80;
wire n_0_0_81;
wire n_0_0_82;
wire n_0_0_83;
wire n_0_0_84;
wire n_0_0_85;
wire n_0_0_86;
wire n_0_0_87;
wire n_0_0_88;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_0_89;
wire n_0_0_90;
wire n_0_0_91;
wire n_0_0_92;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_9;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_40;
wire n_0_0_47;
wire n_0_0_48;
wire n_0_0_49;
wire n_0_0_50;
wire n_0_0_51;
wire n_0_0_52;
wire n_0_0_53;
wire n_0_0_54;
wire n_0_0_55;
wire n_0_0_56;
wire n_0_0_57;
wire n_0_0_58;
wire n_0_0_59;
wire n_0_0_60;
wire n_0_0_61;
wire n_0_0_62;
wire n_0_0_63;
wire n_0_0_64;
wire n_0_0_65;
wire n_0_32;
wire n_0_0_66;
wire n_0_0_67;
wire n_0_33;
wire n_0_0_68;
wire n_0_0_69;
wire n_0_0_70;
wire n_0_0_76;
wire n_0_0_77;
wire n_0_0_78;
wire n_0_0_93;
wire n_0_0_94;


NAND2_X1 i_0_0_155 (.ZN (n_0_0_94), .A1 (\afterB[29] ), .A2 (\afterA[29] ));
INV_X1 i_0_0_154 (.ZN (n_0_0_93), .A (n_0_0_94));
NAND2_X1 i_0_0_153 (.ZN (n_0_0_78), .A1 (\afterB[30] ), .A2 (\afterA[30] ));
AND3_X1 i_0_0_152 (.ZN (n_0_0_77), .A1 (n_0_0_70), .A2 (n_0_0_78), .A3 (n_0_0_94));
NOR2_X1 i_0_0_151 (.ZN (n_0_0_76), .A1 (\afterB[30] ), .A2 (\afterA[30] ));
INV_X1 i_0_0_150 (.ZN (n_0_0_70), .A (n_0_0_76));
NOR4_X1 i_0_0_149 (.ZN (n_0_0_69), .A1 (\afterA[26] ), .A2 (\afterA[23] ), .A3 (\afterA[29] ), .A4 (\afterA[28] ));
NOR4_X1 i_0_0_125 (.ZN (n_0_0_68), .A1 (\afterA[25] ), .A2 (\afterA[24] ), .A3 (\afterA[30] ), .A4 (\afterA[27] ));
NAND2_X1 i_0_0_124 (.ZN (n_0_33), .A1 (n_0_0_69), .A2 (n_0_0_68));
NOR4_X1 i_0_0_123 (.ZN (n_0_0_67), .A1 (\afterB[26] ), .A2 (\afterB[23] ), .A3 (\afterB[29] ), .A4 (\afterB[28] ));
NOR4_X1 i_0_0_122 (.ZN (n_0_0_66), .A1 (\afterB[25] ), .A2 (\afterB[24] ), .A3 (\afterB[30] ), .A4 (\afterB[27] ));
NAND2_X1 i_0_0_121 (.ZN (n_0_32), .A1 (n_0_0_67), .A2 (n_0_0_66));
INV_X1 i_0_0_120 (.ZN (n_0_0_65), .A (\afterB[24] ));
INV_X1 i_0_0_119 (.ZN (n_0_0_64), .A (\afterA[24] ));
NAND2_X1 i_0_0_118 (.ZN (n_0_0_63), .A1 (\afterB[25] ), .A2 (\afterA[25] ));
NAND2_X1 i_0_0_117 (.ZN (n_0_0_62), .A1 (\afterB[26] ), .A2 (\afterA[26] ));
OAI21_X1 i_0_0_116 (.ZN (n_0_0_61), .A (n_0_0_62), .B1 (\afterB[26] ), .B2 (\afterA[26] ));
NOR2_X1 i_0_0_115 (.ZN (n_0_0_60), .A1 (n_0_0_63), .A2 (n_0_0_61));
AOI21_X1 i_0_0_114 (.ZN (n_0_0_59), .A (n_0_0_60), .B1 (n_0_0_63), .B2 (n_0_0_61));
INV_X1 i_0_0_113 (.ZN (n_0_0_58), .A (n_0_0_59));
OAI21_X1 i_0_0_112 (.ZN (n_0_0_57), .A (n_0_0_63), .B1 (\afterB[25] ), .B2 (\afterA[25] ));
NOR3_X1 i_0_0_111 (.ZN (n_0_0_56), .A1 (n_0_0_65), .A2 (n_0_0_64), .A3 (n_0_0_57));
INV_X1 i_0_0_110 (.ZN (n_0_0_55), .A (n_0_0_56));
AOI21_X1 i_0_0_109 (.ZN (n_0_0_54), .A (n_0_0_4), .B1 (n_0_0_9), .B2 (n_0_0_3));
OAI21_X1 i_0_0_108 (.ZN (n_0_0_53), .A (n_0_0_57), .B1 (n_0_0_65), .B2 (n_0_0_64));
AOI21_X1 i_0_0_107 (.ZN (n_0_0_52), .A (n_0_0_56), .B1 (n_0_0_54), .B2 (n_0_0_53));
NOR2_X1 i_0_0_106 (.ZN (n_0_0_51), .A1 (n_0_0_58), .A2 (n_0_0_52));
NOR2_X1 i_0_0_105 (.ZN (n_0_0_50), .A1 (n_0_0_60), .A2 (n_0_0_51));
NAND2_X1 i_0_0_104 (.ZN (n_0_0_49), .A1 (\afterB[27] ), .A2 (\afterA[27] ));
OAI21_X1 i_0_0_103 (.ZN (n_0_0_48), .A (n_0_0_49), .B1 (\afterB[27] ), .B2 (\afterA[27] ));
XNOR2_X1 i_0_0_102 (.ZN (n_0_0_47), .A (n_0_0_62), .B (n_0_0_48));
OAI22_X1 i_0_0_101 (.ZN (n_0_0_40), .A1 (n_0_0_62), .A2 (n_0_0_48), .B1 (n_0_0_50), .B2 (n_0_0_47));
XNOR2_X1 i_0_0_100 (.ZN (n_0_0_21), .A (\afterB[28] ), .B (\afterA[28] ));
XOR2_X1 i_0_0_99 (.Z (n_0_0_20), .A (n_0_0_49), .B (n_0_0_21));
XNOR2_X1 i_0_0_98 (.ZN (n_0_0_19), .A (n_0_0_40), .B (n_0_0_20));
XNOR2_X1 i_0_0_97 (.ZN (n_0_0_18), .A (n_0_0_9), .B (n_0_0_17));
NAND2_X1 i_0_0_96 (.ZN (n_0_0_17), .A1 (n_0_0_16), .A2 (n_0_0_3));
INV_X1 i_0_0_95 (.ZN (n_0_0_16), .A (n_0_0_4));
XNOR2_X1 i_0_0_94 (.ZN (n_0_0_9), .A (\afterB[24] ), .B (\afterA[24] ));
NOR3_X1 i_0_0_93 (.ZN (n_0_0_4), .A1 (\afterB[23] ), .A2 (\MP[47] ), .A3 (\afterA[23] ));
NAND3_X1 i_0_0_92 (.ZN (n_0_0_3), .A1 (\afterB[23] ), .A2 (\MP[47] ), .A3 (\afterA[23] ));
NAND4_X1 i_0_0_91 (.ZN (n_0_0_92), .A1 (\afterB[26] ), .A2 (\afterB[25] ), .A3 (\afterB[24] ), .A4 (\afterB[23] ));
NAND4_X1 i_0_0_90 (.ZN (n_0_0_91), .A1 (\afterB[30] ), .A2 (\afterB[29] ), .A3 (\afterB[28] ), .A4 (\afterB[27] ));
NAND4_X1 i_0_0_89 (.ZN (n_0_0_90), .A1 (\afterA[26] ), .A2 (\afterA[25] ), .A3 (\afterA[24] ), .A4 (\afterA[23] ));
NAND4_X1 i_0_0_88 (.ZN (n_0_0_89), .A1 (\afterA[30] ), .A2 (\afterA[29] ), .A3 (\afterA[28] ), .A4 (\afterA[27] ));
OAI22_X1 i_0_0_87 (.ZN (Exception), .A1 (n_0_0_92), .A2 (n_0_0_91), .B1 (n_0_0_90), .B2 (n_0_0_89));
MUX2_X1 i_0_0_148 (.Z (n_0_57), .A (\MP[45] ), .B (\MP[46] ), .S (\MP[47] ));
MUX2_X1 i_0_0_147 (.Z (n_0_56), .A (\MP[44] ), .B (\MP[45] ), .S (\MP[47] ));
MUX2_X1 i_0_0_146 (.Z (n_0_55), .A (\MP[43] ), .B (\MP[44] ), .S (\MP[47] ));
MUX2_X1 i_0_0_145 (.Z (n_0_54), .A (\MP[42] ), .B (\MP[43] ), .S (\MP[47] ));
MUX2_X1 i_0_0_144 (.Z (n_0_53), .A (\MP[41] ), .B (\MP[42] ), .S (\MP[47] ));
MUX2_X1 i_0_0_143 (.Z (n_0_52), .A (\MP[40] ), .B (\MP[41] ), .S (\MP[47] ));
MUX2_X1 i_0_0_142 (.Z (n_0_51), .A (\MP[39] ), .B (\MP[40] ), .S (\MP[47] ));
MUX2_X1 i_0_0_141 (.Z (n_0_50), .A (\MP[38] ), .B (\MP[39] ), .S (\MP[47] ));
MUX2_X1 i_0_0_140 (.Z (n_0_49), .A (\MP[37] ), .B (\MP[38] ), .S (\MP[47] ));
MUX2_X1 i_0_0_139 (.Z (n_0_48), .A (\MP[36] ), .B (\MP[37] ), .S (\MP[47] ));
MUX2_X1 i_0_0_138 (.Z (n_0_47), .A (\MP[35] ), .B (\MP[36] ), .S (\MP[47] ));
MUX2_X1 i_0_0_137 (.Z (n_0_46), .A (\MP[34] ), .B (\MP[35] ), .S (\MP[47] ));
MUX2_X1 i_0_0_136 (.Z (n_0_45), .A (\MP[33] ), .B (\MP[34] ), .S (\MP[47] ));
MUX2_X1 i_0_0_135 (.Z (n_0_44), .A (\MP[32] ), .B (\MP[33] ), .S (\MP[47] ));
MUX2_X1 i_0_0_134 (.Z (n_0_43), .A (\MP[31] ), .B (\MP[32] ), .S (\MP[47] ));
MUX2_X1 i_0_0_133 (.Z (n_0_42), .A (\MP[30] ), .B (\MP[31] ), .S (\MP[47] ));
MUX2_X1 i_0_0_132 (.Z (n_0_41), .A (\MP[29] ), .B (\MP[30] ), .S (\MP[47] ));
MUX2_X1 i_0_0_131 (.Z (n_0_40), .A (\MP[28] ), .B (\MP[29] ), .S (\MP[47] ));
MUX2_X1 i_0_0_130 (.Z (n_0_39), .A (\MP[27] ), .B (\MP[28] ), .S (\MP[47] ));
MUX2_X1 i_0_0_129 (.Z (n_0_38), .A (\MP[26] ), .B (\MP[27] ), .S (\MP[47] ));
MUX2_X1 i_0_0_128 (.Z (n_0_37), .A (\MP[25] ), .B (\MP[26] ), .S (\MP[47] ));
MUX2_X1 i_0_0_127 (.Z (n_0_36), .A (\MP[24] ), .B (\MP[25] ), .S (\MP[47] ));
MUX2_X1 i_0_0_126 (.Z (n_0_35), .A (\MP[23] ), .B (\MP[24] ), .S (\MP[47] ));
NOR2_X1 i_0_0_86 (.ZN (n_0_0_88), .A1 (\MP[21] ), .A2 (\MP[20] ));
NOR4_X1 i_0_0_85 (.ZN (n_0_0_87), .A1 (\MP[19] ), .A2 (\MP[18] ), .A3 (\MP[17] ), .A4 (\MP[16] ));
NOR4_X1 i_0_0_84 (.ZN (n_0_0_86), .A1 (\MP[11] ), .A2 (\MP[10] ), .A3 (\MP[9] ), .A4 (\MP[8] ));
NOR4_X1 i_0_0_83 (.ZN (n_0_0_85), .A1 (\MP[15] ), .A2 (\MP[14] ), .A3 (\MP[13] ), .A4 (\MP[12] ));
NOR4_X1 i_0_0_82 (.ZN (n_0_0_84), .A1 (\MP[3] ), .A2 (\MP[2] ), .A3 (\MP[1] ), .A4 (\MP[0] ));
NOR4_X1 i_0_0_81 (.ZN (n_0_0_83), .A1 (\MP[7] ), .A2 (\MP[6] ), .A3 (\MP[5] ), .A4 (\MP[4] ));
AND4_X1 i_0_0_80 (.ZN (n_0_0_82), .A1 (n_0_0_86), .A2 (n_0_0_85), .A3 (n_0_0_84), .A4 (n_0_0_83));
NAND3_X1 i_0_0_79 (.ZN (n_0_0_81), .A1 (n_0_0_88), .A2 (n_0_0_87), .A3 (n_0_0_82));
OAI211_X1 i_0_0_78 (.ZN (n_0_0_80), .A (\MP[47] ), .B (\MP[23] ), .C1 (n_0_0_81), .C2 (\MP[22] ));
NAND2_X1 i_0_0_77 (.ZN (n_0_0_79), .A1 (n_0_0_81), .A2 (\MP[22] ));
OAI21_X1 i_0_0_76 (.ZN (n_0_34), .A (n_0_0_80), .B1 (n_0_0_79), .B2 (\MP[47] ));
AOI21_X1 i_0_0_75 (.ZN (n_0_0_75), .A (n_0_0_94), .B1 (n_0_0_70), .B2 (n_0_0_78));
NAND2_X1 i_0_0_74 (.ZN (n_0_0_74), .A1 (\afterB[28] ), .A2 (\afterA[28] ));
NOR2_X1 i_0_0_73 (.ZN (n_0_0_73), .A1 (\afterB[29] ), .A2 (\afterA[29] ));
OAI21_X1 i_0_0_72 (.ZN (n_0_0_72), .A (n_0_0_74), .B1 (n_0_0_73), .B2 (n_0_0_93));
OR3_X1 i_0_0_71 (.ZN (n_0_0_71), .A1 (n_0_0_93), .A2 (n_0_0_73), .A3 (n_0_0_74));
NAND2_X1 i_0_0_70 (.ZN (n_0_0_46), .A1 (n_0_0_40), .A2 (n_0_0_20));
OAI21_X1 i_0_0_69 (.ZN (n_0_0_45), .A (n_0_0_46), .B1 (n_0_0_21), .B2 (n_0_0_49));
NAND2_X1 i_0_0_68 (.ZN (n_0_0_44), .A1 (n_0_0_72), .A2 (n_0_0_45));
AND2_X1 i_0_0_67 (.ZN (n_0_0_43), .A1 (n_0_0_71), .A2 (n_0_0_44));
INV_X1 i_0_0_66 (.ZN (n_0_0_42), .A (n_0_0_43));
NOR2_X1 i_0_0_65 (.ZN (n_0_0_41), .A1 (n_0_0_75), .A2 (n_0_0_42));
NOR3_X1 i_0_0_64 (.ZN (n_0_0_39), .A1 (n_0_0_76), .A2 (n_0_0_41), .A3 (n_0_0_77));
NOR3_X1 i_0_0_63 (.ZN (n_0_0_38), .A1 (n_0_0_42), .A2 (n_0_0_70), .A3 (n_0_0_75));
OR2_X1 i_0_0_62 (.ZN (n_0_0_37), .A1 (n_0_0_75), .A2 (n_0_0_77));
XNOR2_X1 i_0_0_61 (.ZN (n_0_0_36), .A (n_0_0_43), .B (n_0_0_37));
OAI21_X1 i_0_0_60 (.ZN (n_0_0_35), .A (n_0_0_36), .B1 (n_0_0_38), .B2 (n_0_0_39));
NOR4_X1 i_0_0_59 (.ZN (n_0_0_34), .A1 (\MP_final[18] ), .A2 (\MP_final[17] ), .A3 (\MP_final[16] ), .A4 (\MP_final[15] ));
NOR4_X1 i_0_0_58 (.ZN (n_0_0_33), .A1 (\MP_final[22] ), .A2 (\MP_final[21] ), .A3 (\MP_final[20] ), .A4 (\MP_final[19] ));
NAND2_X1 i_0_0_57 (.ZN (n_0_0_32), .A1 (n_0_0_34), .A2 (n_0_0_33));
NOR4_X1 i_0_0_56 (.ZN (n_0_0_31), .A1 (\MP_final[10] ), .A2 (\MP_final[9] ), .A3 (\MP_final[8] ), .A4 (\MP_final[7] ));
NOR4_X1 i_0_0_55 (.ZN (n_0_0_30), .A1 (\MP_final[14] ), .A2 (\MP_final[13] ), .A3 (\MP_final[12] ), .A4 (\MP_final[11] ));
NOR3_X1 i_0_0_54 (.ZN (n_0_0_29), .A1 (\MP_final[5] ), .A2 (\MP_final[4] ), .A3 (\MP_final[1] ));
NOR4_X1 i_0_0_53 (.ZN (n_0_0_28), .A1 (\MP_final[6] ), .A2 (\MP_final[3] ), .A3 (\MP_final[2] ), .A4 (\MP_final[0] ));
NAND4_X1 i_0_0_52 (.ZN (n_0_0_27), .A1 (n_0_0_31), .A2 (n_0_0_30), .A3 (n_0_0_29), .A4 (n_0_0_28));
NOR2_X1 i_0_0_51 (.ZN (n_0_0_26), .A1 (n_0_0_32), .A2 (n_0_0_27));
INV_X1 i_0_0_50 (.ZN (n_0_0_25), .A (n_0_0_26));
NOR2_X1 i_0_0_49 (.ZN (n_0_0_24), .A1 (Exception), .A2 (n_0_0_25));
NOR2_X1 i_0_0_48 (.ZN (Overflow), .A1 (n_0_0_35), .A2 (n_0_0_24));
NOR3_X1 i_0_0_47 (.ZN (n_0_0_23), .A1 (n_0_0_78), .A2 (n_0_0_74), .A3 (n_0_0_46));
AOI21_X1 i_0_0_46 (.ZN (n_0_0_22), .A (n_0_0_38), .B1 (n_0_0_23), .B2 (n_0_0_93));
NOR2_X1 i_0_0_45 (.ZN (Underflow), .A1 (n_0_0_24), .A2 (n_0_0_22));
XNOR2_X1 i_0_0_44 (.ZN (n_0_0_15), .A (\afterB[31] ), .B (\afterA[31] ));
NOR2_X1 i_0_0_43 (.ZN (n_0_31), .A1 (Exception), .A2 (n_0_0_15));
OR2_X1 i_0_0_42 (.ZN (n_0_0_14), .A1 (n_0_0_26), .A2 (Exception));
OR2_X1 i_0_0_41 (.ZN (n_0_0_13), .A1 (n_0_0_35), .A2 (n_0_0_14));
OR2_X1 i_0_0_40 (.ZN (n_0_0_12), .A1 (n_0_0_38), .A2 (n_0_0_14));
OAI21_X1 i_0_0_39 (.ZN (n_0_30), .A (n_0_0_13), .B1 (n_0_0_12), .B2 (n_0_0_36));
AND2_X1 i_0_0_38 (.ZN (n_0_0_11), .A1 (n_0_0_72), .A2 (n_0_0_71));
XNOR2_X1 i_0_0_37 (.ZN (n_0_0_10), .A (n_0_0_45), .B (n_0_0_11));
OAI21_X1 i_0_0_36 (.ZN (n_0_29), .A (n_0_0_13), .B1 (n_0_0_12), .B2 (n_0_0_10));
OAI21_X1 i_0_0_35 (.ZN (n_0_28), .A (n_0_0_13), .B1 (n_0_0_12), .B2 (n_0_0_19));
XNOR2_X1 i_0_0_34 (.ZN (n_0_0_8), .A (n_0_0_50), .B (n_0_0_47));
OAI21_X1 i_0_0_33 (.ZN (n_0_27), .A (n_0_0_13), .B1 (n_0_0_12), .B2 (n_0_0_8));
AND2_X1 i_0_0_32 (.ZN (n_0_0_7), .A1 (n_0_0_58), .A2 (n_0_0_52));
OAI33_X1 i_0_0_31 (.ZN (n_0_26), .A1 (Exception), .A2 (n_0_0_35), .A3 (n_0_0_26), .B1 (n_0_0_12)
    , .B2 (n_0_0_7), .B3 (n_0_0_51));
NAND2_X1 i_0_0_30 (.ZN (n_0_0_6), .A1 (n_0_0_53), .A2 (n_0_0_55));
XOR2_X1 i_0_0_29 (.Z (n_0_0_5), .A (n_0_0_54), .B (n_0_0_6));
OAI21_X1 i_0_0_28 (.ZN (n_0_25), .A (n_0_0_13), .B1 (n_0_0_12), .B2 (n_0_0_5));
OAI21_X1 i_0_0_27 (.ZN (n_0_24), .A (n_0_0_13), .B1 (n_0_0_12), .B2 (n_0_0_18));
XNOR2_X1 i_0_0_26 (.ZN (n_0_0_2), .A (\MP[47] ), .B (\afterA[23] ));
XNOR2_X1 i_0_0_25 (.ZN (n_0_0_1), .A (\afterB[23] ), .B (n_0_0_2));
OAI21_X1 i_0_0_24 (.ZN (n_0_23), .A (n_0_0_13), .B1 (n_0_0_12), .B2 (n_0_0_1));
NOR2_X2 i_0_0_23 (.ZN (n_0_0_0), .A1 (n_0_0_39), .A2 (n_0_0_12));
AND2_X1 i_0_0_22 (.ZN (n_0_22), .A1 (\MP_final[22] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_21 (.ZN (n_0_21), .A1 (\MP_final[21] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_20 (.ZN (n_0_20), .A1 (\MP_final[20] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_19 (.ZN (n_0_19), .A1 (\MP_final[19] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_18 (.ZN (n_0_18), .A1 (\MP_final[18] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_17 (.ZN (n_0_17), .A1 (\MP_final[17] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_16 (.ZN (n_0_16), .A1 (\MP_final[16] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_15 (.ZN (n_0_15), .A1 (\MP_final[15] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_14 (.ZN (n_0_14), .A1 (\MP_final[14] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_13 (.ZN (n_0_13), .A1 (\MP_final[13] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_12 (.ZN (n_0_12), .A1 (\MP_final[12] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_11 (.ZN (n_0_11), .A1 (\MP_final[11] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_10 (.ZN (n_0_10), .A1 (\MP_final[10] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_9 (.ZN (n_0_9), .A1 (\MP_final[9] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_8 (.ZN (n_0_8), .A1 (\MP_final[8] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_7 (.ZN (n_0_7), .A1 (\MP_final[7] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_6 (.ZN (n_0_6), .A1 (\MP_final[6] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_5 (.ZN (n_0_5), .A1 (\MP_final[5] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_4 (.ZN (n_0_4), .A1 (\MP_final[4] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_3 (.ZN (n_0_3), .A1 (\MP_final[3] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_2 (.ZN (n_0_2), .A1 (\MP_final[2] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_1 (.ZN (n_0_1), .A1 (\MP_final[1] ), .A2 (n_0_0_0));
AND2_X1 i_0_0_0 (.ZN (n_0_0), .A1 (\MP_final[0] ), .A2 (n_0_0_0));
datapath__0_4 i_0_6 (.MP_final ({\MP_final[22] , \MP_final[21] , \MP_final[20] , 
    \MP_final[19] , \MP_final[18] , \MP_final[17] , \MP_final[16] , \MP_final[15] , 
    \MP_final[14] , \MP_final[13] , \MP_final[12] , \MP_final[11] , \MP_final[10] , 
    \MP_final[9] , \MP_final[8] , \MP_final[7] , \MP_final[6] , \MP_final[5] , \MP_final[4] , 
    \MP_final[3] , \MP_final[2] , \MP_final[1] , \MP_final[0] }), .p_0 ({1'b0 , 1'b0 , 
    1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 
    1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , n_0_34}), .p_1 ({
    n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, 
    n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, 
    n_0_37, n_0_36, n_0_35}));
Reg regOut (.out ({Out[31], Out[30], Out[29], Out[28], Out[27], Out[26], Out[25], 
    Out[24], Out[23], Out[22], Out[21], Out[20], Out[19], Out[18], Out[17], Out[16], 
    Out[15], Out[14], Out[13], Out[12], Out[11], Out[10], Out[9], Out[8], Out[7], 
    Out[6], Out[5], Out[4], Out[3], Out[2], Out[1], Out[0]}), .clk (clk), .in ({n_0_31, 
    n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, 
    n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, 
    n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0}));
N_Bit_Mult mantissa_multiplier (.Out ({\MP[47] , \MP[46] , \MP[45] , \MP[44] , \MP[43] , 
    \MP[42] , \MP[41] , \MP[40] , \MP[39] , \MP[38] , \MP[37] , \MP[36] , \MP[35] , 
    \MP[34] , \MP[33] , \MP[32] , \MP[31] , \MP[30] , \MP[29] , \MP[28] , \MP[27] , 
    \MP[26] , \MP[25] , \MP[24] , \MP[23] , \MP[22] , \MP[21] , \MP[20] , \MP[19] , 
    \MP[18] , \MP[17] , \MP[16] , \MP[15] , \MP[14] , \MP[13] , \MP[12] , \MP[11] , 
    \MP[10] , \MP[9] , \MP[8] , \MP[7] , \MP[6] , \MP[5] , \MP[4] , \MP[3] , \MP[2] , 
    \MP[1] , \MP[0] }), .A ({n_0_33, \afterA[22] , \afterA[21] , \afterA[20] , \afterA[19] , 
    \afterA[18] , \afterA[17] , \afterA[16] , \afterA[15] , \afterA[14] , \afterA[13] , 
    \afterA[12] , \afterA[11] , \afterA[10] , \afterA[9] , \afterA[8] , \afterA[7] , 
    \afterA[6] , \afterA[5] , \afterA[4] , \afterA[3] , \afterA[2] , \afterA[1] , 
    \afterA[0] }), .B ({n_0_32, \afterB[22] , \afterB[21] , \afterB[20] , \afterB[19] , 
    \afterB[18] , \afterB[17] , \afterB[16] , \afterB[15] , \afterB[14] , \afterB[13] , 
    \afterB[12] , \afterB[11] , \afterB[10] , \afterB[9] , \afterB[8] , \afterB[7] , 
    \afterB[6] , \afterB[5] , \afterB[4] , \afterB[3] , \afterB[2] , \afterB[1] , 
    \afterB[0] }));
Reg__0_18 regA (.out ({\afterA[31] , \afterA[30] , \afterA[29] , \afterA[28] , \afterA[27] , 
    \afterA[26] , \afterA[25] , \afterA[24] , \afterA[23] , \afterA[22] , \afterA[21] , 
    \afterA[20] , \afterA[19] , \afterA[18] , \afterA[17] , \afterA[16] , \afterA[15] , 
    \afterA[14] , \afterA[13] , \afterA[12] , \afterA[11] , \afterA[10] , \afterA[9] , 
    \afterA[8] , \afterA[7] , \afterA[6] , \afterA[5] , \afterA[4] , \afterA[3] , 
    \afterA[2] , \afterA[1] , \afterA[0] }), .clk (clk), .in ({A[31], A[30], A[29], 
    A[28], A[27], A[26], A[25], A[24], A[23], A[22], A[21], A[20], A[19], A[18], 
    A[17], A[16], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], 
    A[5], A[4], A[3], A[2], A[1], A[0]}));
Reg__0_17 regB (.out ({\afterB[31] , \afterB[30] , \afterB[29] , \afterB[28] , \afterB[27] , 
    \afterB[26] , \afterB[25] , \afterB[24] , \afterB[23] , \afterB[22] , \afterB[21] , 
    \afterB[20] , \afterB[19] , \afterB[18] , \afterB[17] , \afterB[16] , \afterB[15] , 
    \afterB[14] , \afterB[13] , \afterB[12] , \afterB[11] , \afterB[10] , \afterB[9] , 
    \afterB[8] , \afterB[7] , \afterB[6] , \afterB[5] , \afterB[4] , \afterB[3] , 
    \afterB[2] , \afterB[1] , \afterB[0] }), .clk (clk), .in ({B[31], B[30], B[29], 
    B[28], B[27], B[26], B[25], B[24], B[23], B[22], B[21], B[20], B[19], B[18], 
    B[17], B[16], B[15], B[14], B[13], B[12], B[11], B[10], B[9], B[8], B[7], B[6], 
    B[5], B[4], B[3], B[2], B[1], B[0]}));

endmodule //float_mult


