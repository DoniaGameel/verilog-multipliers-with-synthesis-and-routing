/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sun Jan  1 16:46:23 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3428632784 */

module datapath(inputB, inputA, result);
   input [31:0]inputB;
   input [31:0]inputA;
   output [63:0]result;

   HA_X1 i_1052 (.A(n_1030), .B(n_1045), .CO(n_1053), .S(n_1052));
   HA_X1 i_1067 (.A(n_1040), .B(n_1046), .CO(n_1069), .S(n_1068));
   HA_X1 i_1071 (.A(n_1056), .B(n_1053), .CO(n_1074), .S(n_1073));
   HA_X1 i_1094 (.A(n_1084), .B(n_1077), .CO(n_1098), .S(n_1097));
   HA_X1 i_1098 (.A(n_1074), .B(n_1072), .CO(n_1103), .S(n_1102));
   HA_X1 i_1121 (.A(n_1078), .B(n_1092), .CO(n_1127), .S(n_1126));
   HA_X1 i_1125 (.A(n_1113), .B(n_1106), .CO(n_1132), .S(n_1131));
   HA_X1 i_1129 (.A(n_1128), .B(n_1101), .CO(n_1137), .S(n_1136));
   HA_X1 i_1151 (.A(n_1114), .B(n_1107), .CO(n_1160), .S(n_1159));
   HA_X1 i_1155 (.A(n_1154), .B(n_1147), .CO(n_1165), .S(n_1164));
   HA_X1 i_1159 (.A(n_1161), .B(n_1130), .CO(n_1170), .S(n_1169));
   HA_X1 i_1163 (.A(n_1135), .B(n_1166), .CO(n_1175), .S(n_1174));
   HA_X1 i_1193 (.A(n_1141), .B(n_1192), .CO(n_1206), .S(n_1205));
   HA_X1 i_1197 (.A(n_1178), .B(n_1163), .CO(n_1211), .S(n_1210));
   HA_X1 i_1201 (.A(n_1168), .B(n_1207), .CO(n_1216), .S(n_1215));
   HA_X1 i_1205 (.A(n_1175), .B(n_1173), .CO(n_1221), .S(n_1220));
   HA_X1 i_1235 (.A(n_1186), .B(n_1179), .CO(n_1252), .S(n_1251));
   HA_X1 i_1239 (.A(n_1244), .B(n_1238), .CO(n_1257), .S(n_1256));
   HA_X1 i_1243 (.A(n_1224), .B(n_1253), .CO(n_1262), .S(n_1261));
   HA_X1 i_1247 (.A(n_1214), .B(n_1258), .CO(n_1267), .S(n_1266));
   HA_X1 i_1251 (.A(n_1221), .B(n_1219), .CO(n_1272), .S(n_1271));
   HA_X1 i_1280 (.A(n_1239), .B(n_1232), .CO(n_1302), .S(n_1301));
   HA_X1 i_1284 (.A(n_1245), .B(n_1296), .CO(n_1307), .S(n_1306));
   HA_X1 i_1288 (.A(n_1282), .B(n_1275), .CO(n_1312), .S(n_1311));
   HA_X1 i_1292 (.A(n_1303), .B(n_1260), .CO(n_1317), .S(n_1316));
   HA_X1 i_1296 (.A(n_1313), .B(n_1308), .CO(n_1322), .S(n_1321));
   HA_X1 i_1300 (.A(n_1272), .B(n_1270), .CO(n_1327), .S(n_1326));
   HA_X1 i_1337 (.A(n_1283), .B(n_1276), .CO(n_1365), .S(n_1364));
   HA_X1 i_1341 (.A(n_1351), .B(n_1344), .CO(n_1370), .S(n_1369));
   HA_X1 i_1345 (.A(n_1330), .B(n_1366), .CO(n_1375), .S(n_1374));
   HA_X1 i_1349 (.A(n_1310), .B(n_1315), .CO(n_1380), .S(n_1379));
   HA_X1 i_1353 (.A(n_1320), .B(n_1376), .CO(n_1385), .S(n_1384));
   HA_X1 i_1357 (.A(n_1325), .B(n_1327), .CO(n_1390), .S(n_1389));
   HA_X1 i_1394 (.A(n_1345), .B(n_1338), .CO(n_1428), .S(n_1427));
   HA_X1 i_1398 (.A(n_1359), .B(n_1420), .CO(n_1433), .S(n_1432));
   HA_X1 i_1402 (.A(n_1407), .B(n_1400), .CO(n_1438), .S(n_1437));
   HA_X1 i_1406 (.A(n_1368), .B(n_1429), .CO(n_1443), .S(n_1442));
   HA_X1 i_1410 (.A(n_1378), .B(n_1439), .CO(n_1448), .S(n_1447));
   HA_X1 i_1414 (.A(n_1444), .B(n_1383), .CO(n_1453), .S(n_1452));
   HA_X1 i_1418 (.A(n_1449), .B(n_1390), .CO(n_1458), .S(n_1457));
   HA_X1 i_1454 (.A(n_1415), .B(n_1408), .CO(n_1495), .S(n_1494));
   HA_X1 i_1458 (.A(n_1394), .B(n_1431), .CO(n_1500), .S(n_1499));
   HA_X1 i_1462 (.A(n_1489), .B(n_1482), .CO(n_1505), .S(n_1504));
   HA_X1 i_1466 (.A(n_1468), .B(n_1461), .CO(n_1510), .S(n_1509));
   HA_X1 i_1470 (.A(n_1441), .B(n_1436), .CO(n_1515), .S(n_1514));
   HA_X1 i_1474 (.A(n_1446), .B(n_1511), .CO(n_1520), .S(n_1519));
   HA_X1 i_1478 (.A(n_1516), .B(n_1451), .CO(n_1525), .S(n_1524));
   HA_X1 i_1482 (.A(n_1456), .B(n_1458), .CO(n_1530), .S(n_1529));
   HA_X1 i_1526 (.A(n_1476), .B(n_1469), .CO(n_1575), .S(n_1574));
   HA_X1 i_1530 (.A(n_1498), .B(n_1561), .CO(n_1580), .S(n_1579));
   HA_X1 i_1534 (.A(n_1547), .B(n_1540), .CO(n_1585), .S(n_1584));
   HA_X1 i_1538 (.A(n_1503), .B(n_1576), .CO(n_1590), .S(n_1589));
   HA_X1 i_1542 (.A(n_1508), .B(n_1513), .CO(n_1595), .S(n_1594));
   HA_X1 i_1546 (.A(n_1581), .B(n_1518), .CO(n_1600), .S(n_1599));
   HA_X1 i_1550 (.A(n_1523), .B(n_1596), .CO(n_1605), .S(n_1604));
   HA_X1 i_1554 (.A(n_1528), .B(n_1530), .CO(n_1610), .S(n_1609));
   HA_X1 i_1598 (.A(n_1555), .B(n_1548), .CO(n_1655), .S(n_1654));
   HA_X1 i_1602 (.A(n_1534), .B(n_1578), .CO(n_1660), .S(n_1659));
   HA_X1 i_1606 (.A(n_1647), .B(n_1641), .CO(n_1665), .S(n_1664));
   HA_X1 i_1610 (.A(n_1627), .B(n_1620), .CO(n_1670), .S(n_1669));
   HA_X1 i_1614 (.A(n_1656), .B(n_1588), .CO(n_1675), .S(n_1674));
   HA_X1 i_1618 (.A(n_1661), .B(n_1593), .CO(n_1680), .S(n_1679));
   HA_X1 i_1622 (.A(n_1666), .B(n_1676), .CO(n_1685), .S(n_1684));
   HA_X1 i_1626 (.A(n_1681), .B(n_1603), .CO(n_1690), .S(n_1689));
   HA_X1 i_1630 (.A(n_1608), .B(n_1610), .CO(n_1695), .S(n_1694));
   HA_X1 i_1673 (.A(n_1642), .B(n_1635), .CO(n_1739), .S(n_1738));
   HA_X1 i_1677 (.A(n_1621), .B(n_1614), .CO(n_1744), .S(n_1743));
   HA_X1 i_1681 (.A(n_1648), .B(n_1733), .CO(n_1749), .S(n_1748));
   HA_X1 i_1685 (.A(n_1719), .B(n_1712), .CO(n_1754), .S(n_1753));
   HA_X1 i_1689 (.A(n_1698), .B(n_1663), .CO(n_1759), .S(n_1758));
   HA_X1 i_1693 (.A(n_1740), .B(n_1673), .CO(n_1764), .S(n_1763));
   HA_X1 i_1697 (.A(n_1678), .B(n_1755), .CO(n_1769), .S(n_1768));
   HA_X1 i_1701 (.A(n_1760), .B(n_1765), .CO(n_1774), .S(n_1773));
   HA_X1 i_1705 (.A(n_1688), .B(n_1770), .CO(n_1779), .S(n_1778));
   HA_X1 i_1709 (.A(n_1693), .B(n_1695), .CO(n_1784), .S(n_1783));
   HA_X1 i_1760 (.A(n_1720), .B(n_1713), .CO(n_1836), .S(n_1835));
   HA_X1 i_1764 (.A(n_1699), .B(n_1742), .CO(n_1841), .S(n_1840));
   HA_X1 i_1768 (.A(n_1815), .B(n_1808), .CO(n_1846), .S(n_1845));
   HA_X1 i_1772 (.A(n_1794), .B(n_1787), .CO(n_1851), .S(n_1850));
   HA_X1 i_1776 (.A(n_1837), .B(n_1829), .CO(n_1856), .S(n_1855));
   HA_X1 i_1780 (.A(n_1752), .B(n_1842), .CO(n_1861), .S(n_1860));
   HA_X1 i_1784 (.A(n_1762), .B(n_1852), .CO(n_1866), .S(n_1865));
   HA_X1 i_1788 (.A(n_1857), .B(n_1772), .CO(n_1871), .S(n_1870));
   HA_X1 i_1792 (.A(n_1777), .B(n_1867), .CO(n_1876), .S(n_1875));
   HA_X1 i_1796 (.A(n_1782), .B(n_1877), .CO(n_1881), .S(n_1880));
   HA_X1 i_1847 (.A(n_1816), .B(n_1809), .CO(n_1933), .S(n_1932));
   HA_X1 i_1851 (.A(n_1795), .B(n_1788), .CO(n_1938), .S(n_1937));
   HA_X1 i_1855 (.A(n_1830), .B(n_1925), .CO(n_1943), .S(n_1942));
   HA_X1 i_1859 (.A(n_1912), .B(n_1905), .CO(n_1948), .S(n_1947));
   HA_X1 i_1863 (.A(n_1891), .B(n_1884), .CO(n_1953), .S(n_1952));
   HA_X1 i_1867 (.A(n_1934), .B(n_1849), .CO(n_1958), .S(n_1957));
   HA_X1 i_1871 (.A(n_1854), .B(n_1859), .CO(n_1963), .S(n_1962));
   HA_X1 i_1875 (.A(n_1949), .B(n_1944), .CO(n_1968), .S(n_1967));
   HA_X1 i_1879 (.A(n_1959), .B(n_1869), .CO(n_1973), .S(n_1972));
   HA_X1 i_1883 (.A(n_1969), .B(n_1874), .CO(n_1978), .S(n_1977));
   HA_X1 i_1887 (.A(n_1879), .B(n_1979), .CO(n_1983), .S(n_1982));
   HA_X1 i_1937 (.A(n_1920), .B(n_1913), .CO(n_2034), .S(n_2033));
   HA_X1 i_1941 (.A(n_1899), .B(n_1892), .CO(n_2039), .S(n_2038));
   HA_X1 i_1945 (.A(n_1936), .B(n_1926), .CO(n_2044), .S(n_2043));
   HA_X1 i_1949 (.A(n_2021), .B(n_2014), .CO(n_2049), .S(n_2048));
   HA_X1 i_1953 (.A(n_2000), .B(n_1993), .CO(n_2054), .S(n_2053));
   HA_X1 i_1957 (.A(n_1941), .B(n_2040), .CO(n_2059), .S(n_2058));
   HA_X1 i_1961 (.A(n_1951), .B(n_1946), .CO(n_2064), .S(n_2063));
   HA_X1 i_1965 (.A(n_1961), .B(n_1956), .CO(n_2069), .S(n_2068));
   HA_X1 i_1969 (.A(n_2050), .B(n_2065), .CO(n_2074), .S(n_2073));
   HA_X1 i_1973 (.A(n_1966), .B(n_1971), .CO(n_2079), .S(n_2078));
   HA_X1 i_1977 (.A(n_1976), .B(n_2075), .CO(n_2084), .S(n_2083));
   HA_X1 i_1981 (.A(n_1981), .B(n_1983), .CO(n_2089), .S(n_2088));
   HA_X1 i_2039 (.A(n_2015), .B(n_2008), .CO(n_2148), .S(n_2147));
   HA_X1 i_2043 (.A(n_1994), .B(n_1987), .CO(n_2153), .S(n_2152));
   HA_X1 i_2047 (.A(n_2037), .B(n_2134), .CO(n_2158), .S(n_2157));
   HA_X1 i_2051 (.A(n_2120), .B(n_2113), .CO(n_2163), .S(n_2162));
   HA_X1 i_2055 (.A(n_2099), .B(n_2092), .CO(n_2168), .S(n_2167));
   HA_X1 i_2059 (.A(n_2149), .B(n_2141), .CO(n_2173), .S(n_2172));
   HA_X1 i_2063 (.A(n_2052), .B(n_2047), .CO(n_2178), .S(n_2177));
   HA_X1 i_2067 (.A(n_2169), .B(n_2164), .CO(n_2183), .S(n_2182));
   HA_X1 i_2071 (.A(n_2067), .B(n_2179), .CO(n_2188), .S(n_2187));
   HA_X1 i_2075 (.A(n_2072), .B(n_2077), .CO(n_2193), .S(n_2192));
   HA_X1 i_2079 (.A(n_2082), .B(n_2189), .CO(n_2198), .S(n_2197));
   HA_X1 i_2083 (.A(n_2087), .B(n_2199), .CO(n_2203), .S(n_2202));
   HA_X1 i_2141 (.A(n_2128), .B(n_2121), .CO(n_2262), .S(n_2261));
   HA_X1 i_2145 (.A(n_2107), .B(n_2100), .CO(n_2267), .S(n_2266));
   HA_X1 i_2149 (.A(n_2151), .B(n_2142), .CO(n_2272), .S(n_2271));
   HA_X1 i_2153 (.A(n_2248), .B(n_2241), .CO(n_2277), .S(n_2276));
   HA_X1 i_2157 (.A(n_2227), .B(n_2220), .CO(n_2282), .S(n_2281));
   HA_X1 i_2161 (.A(n_2206), .B(n_2156), .CO(n_2287), .S(n_2286));
   HA_X1 i_2165 (.A(n_2263), .B(n_2166), .CO(n_2292), .S(n_2291));
   HA_X1 i_2169 (.A(n_2273), .B(n_2176), .CO(n_2297), .S(n_2296));
   HA_X1 i_2173 (.A(n_2283), .B(n_2278), .CO(n_2302), .S(n_2301));
   HA_X1 i_2177 (.A(n_2181), .B(n_2293), .CO(n_2307), .S(n_2306));
   HA_X1 i_2181 (.A(n_2298), .B(n_2191), .CO(n_2312), .S(n_2311));
   HA_X1 i_2185 (.A(n_2308), .B(n_2196), .CO(n_2317), .S(n_2316));
   HA_X1 i_2189 (.A(n_2201), .B(n_2318), .CO(n_2322), .S(n_2321));
   HA_X1 i_2246 (.A(n_2249), .B(n_2242), .CO(n_2380), .S(n_2379));
   HA_X1 i_2250 (.A(n_2228), .B(n_2221), .CO(n_2385), .S(n_2384));
   HA_X1 i_2254 (.A(n_2207), .B(n_2270), .CO(n_2390), .S(n_2389));
   HA_X1 i_2258 (.A(n_2255), .B(n_2374), .CO(n_2395), .S(n_2394));
   HA_X1 i_2262 (.A(n_2360), .B(n_2353), .CO(n_2400), .S(n_2399));
   HA_X1 i_2266 (.A(n_2339), .B(n_2332), .CO(n_2405), .S(n_2404));
   HA_X1 i_2270 (.A(n_2386), .B(n_2381), .CO(n_2410), .S(n_2409));
   HA_X1 i_2274 (.A(n_2280), .B(n_2275), .CO(n_2415), .S(n_2414));
   HA_X1 i_2278 (.A(n_2295), .B(n_2290), .CO(n_2420), .S(n_2419));
   HA_X1 i_2282 (.A(n_2401), .B(n_2396), .CO(n_2425), .S(n_2424));
   HA_X1 i_2286 (.A(n_2416), .B(n_2411), .CO(n_2430), .S(n_2429));
   HA_X1 i_2290 (.A(n_2421), .B(n_2310), .CO(n_2435), .S(n_2434));
   HA_X1 i_2294 (.A(n_2431), .B(n_2315), .CO(n_2440), .S(n_2439));
   HA_X1 i_2298 (.A(n_2320), .B(n_2441), .CO(n_2445), .S(n_2444));
   HA_X1 i_2363 (.A(n_2361), .B(n_2354), .CO(n_2511), .S(n_2510));
   HA_X1 i_2367 (.A(n_2340), .B(n_2333), .CO(n_2516), .S(n_2515));
   HA_X1 i_2371 (.A(n_2388), .B(n_2383), .CO(n_2521), .S(n_2520));
   HA_X1 i_2375 (.A(n_2490), .B(n_2483), .CO(n_2526), .S(n_2525));
   HA_X1 i_2379 (.A(n_2469), .B(n_2462), .CO(n_2531), .S(n_2530));
   HA_X1 i_2383 (.A(n_2448), .B(n_2393), .CO(n_2536), .S(n_2535));
   HA_X1 i_2387 (.A(n_2512), .B(n_2504), .CO(n_2541), .S(n_2540));
   HA_X1 i_2391 (.A(n_2403), .B(n_2398), .CO(n_2546), .S(n_2545));
   HA_X1 i_2395 (.A(n_2413), .B(n_2532), .CO(n_2551), .S(n_2550));
   HA_X1 i_2399 (.A(n_2537), .B(n_2418), .CO(n_2556), .S(n_2555));
   HA_X1 i_2403 (.A(n_2542), .B(n_2423), .CO(n_2561), .S(n_2560));
   HA_X1 i_2407 (.A(n_2433), .B(n_2552), .CO(n_2566), .S(n_2565));
   HA_X1 i_2411 (.A(n_2562), .B(n_2438), .CO(n_2571), .S(n_2570));
   HA_X1 i_2415 (.A(n_2443), .B(n_2572), .CO(n_2576), .S(n_2575));
   HA_X1 i_2480 (.A(n_2491), .B(n_2484), .CO(n_2642), .S(n_2641));
   HA_X1 i_2484 (.A(n_2470), .B(n_2463), .CO(n_2647), .S(n_2646));
   HA_X1 i_2488 (.A(n_2449), .B(n_2519), .CO(n_2652), .S(n_2651));
   HA_X1 i_2492 (.A(n_2505), .B(n_2634), .CO(n_2657), .S(n_2656));
   HA_X1 i_2496 (.A(n_2621), .B(n_2614), .CO(n_2662), .S(n_2661));
   HA_X1 i_2500 (.A(n_2600), .B(n_2593), .CO(n_2667), .S(n_2666));
   HA_X1 i_2504 (.A(n_2579), .B(n_2648), .CO(n_2672), .S(n_2671));
   HA_X1 i_2508 (.A(n_2534), .B(n_2529), .CO(n_2677), .S(n_2676));
   HA_X1 i_2512 (.A(n_2653), .B(n_2544), .CO(n_2682), .S(n_2681));
   HA_X1 i_2516 (.A(n_2668), .B(n_2663), .CO(n_2687), .S(n_2686));
   HA_X1 i_2520 (.A(n_2549), .B(n_2678), .CO(n_2692), .S(n_2691));
   HA_X1 i_2524 (.A(n_2554), .B(n_2683), .CO(n_2697), .S(n_2696));
   HA_X1 i_2528 (.A(n_2564), .B(n_2688), .CO(n_2702), .S(n_2701));
   HA_X1 i_2532 (.A(n_2569), .B(n_2698), .CO(n_2707), .S(n_2706));
   HA_X1 i_2536 (.A(n_2574), .B(n_2576), .CO(n_2712), .S(n_2711));
   HA_X1 i_2600 (.A(n_2629), .B(n_2622), .CO(n_2777), .S(n_2776));
   HA_X1 i_2604 (.A(n_2608), .B(n_2601), .CO(n_2782), .S(n_2781));
   HA_X1 i_2608 (.A(n_2587), .B(n_2580), .CO(n_2787), .S(n_2786));
   HA_X1 i_2612 (.A(n_2645), .B(n_2635), .CO(n_2792), .S(n_2791));
   HA_X1 i_2616 (.A(n_2764), .B(n_2757), .CO(n_2797), .S(n_2796));
   HA_X1 i_2620 (.A(n_2743), .B(n_2736), .CO(n_2802), .S(n_2801));
   HA_X1 i_2624 (.A(n_2722), .B(n_2715), .CO(n_2807), .S(n_2806));
   HA_X1 i_2628 (.A(n_2788), .B(n_2783), .CO(n_2812), .S(n_2811));
   HA_X1 i_2632 (.A(n_2670), .B(n_2665), .CO(n_2817), .S(n_2816));
   HA_X1 i_2636 (.A(n_2793), .B(n_2680), .CO(n_2822), .S(n_2821));
   HA_X1 i_2640 (.A(n_2808), .B(n_2803), .CO(n_2827), .S(n_2826));
   HA_X1 i_2644 (.A(n_2685), .B(n_2818), .CO(n_2832), .S(n_2831));
   HA_X1 i_2648 (.A(n_2690), .B(n_2823), .CO(n_2837), .S(n_2836));
   HA_X1 i_2652 (.A(n_2828), .B(n_2700), .CO(n_2842), .S(n_2841));
   HA_X1 i_2656 (.A(n_2838), .B(n_2705), .CO(n_2847), .S(n_2846));
   HA_X1 i_2660 (.A(n_2710), .B(n_2848), .CO(n_2852), .S(n_2851));
   HA_X1 i_2732 (.A(n_2758), .B(n_2751), .CO(n_2925), .S(n_2924));
   HA_X1 i_2736 (.A(n_2737), .B(n_2730), .CO(n_2930), .S(n_2929));
   HA_X1 i_2740 (.A(n_2716), .B(n_2785), .CO(n_2935), .S(n_2934));
   HA_X1 i_2744 (.A(n_2911), .B(n_2904), .CO(n_2940), .S(n_2939));
   HA_X1 i_2748 (.A(n_2890), .B(n_2883), .CO(n_2945), .S(n_2944));
   HA_X1 i_2752 (.A(n_2869), .B(n_2862), .CO(n_2950), .S(n_2949));
   HA_X1 i_2756 (.A(n_2790), .B(n_2931), .CO(n_2955), .S(n_2954));
   HA_X1 i_2760 (.A(n_2918), .B(n_2805), .CO(n_2960), .S(n_2959));
   HA_X1 i_2764 (.A(n_2795), .B(n_2810), .CO(n_2965), .S(n_2964));
   HA_X1 i_2768 (.A(n_2820), .B(n_2815), .CO(n_2970), .S(n_2969));
   HA_X1 i_2772 (.A(n_2946), .B(n_2941), .CO(n_2975), .S(n_2974));
   HA_X1 i_2776 (.A(n_2961), .B(n_2956), .CO(n_2980), .S(n_2979));
   HA_X1 i_2780 (.A(n_2966), .B(n_2971), .CO(n_2985), .S(n_2984));
   HA_X1 i_2784 (.A(n_2976), .B(n_2840), .CO(n_2990), .S(n_2989));
   HA_X1 i_2788 (.A(n_2986), .B(n_2845), .CO(n_2995), .S(n_2994));
   HA_X1 i_2792 (.A(n_2850), .B(n_2996), .CO(n_3000), .S(n_2999));
   HA_X1 i_2864 (.A(n_2905), .B(n_2898), .CO(n_3073), .S(n_3072));
   HA_X1 i_2868 (.A(n_2884), .B(n_2877), .CO(n_3078), .S(n_3077));
   HA_X1 i_2872 (.A(n_2863), .B(n_2856), .CO(n_3083), .S(n_3082));
   HA_X1 i_2876 (.A(n_2928), .B(n_2919), .CO(n_3088), .S(n_3087));
   HA_X1 i_2880 (.A(n_3059), .B(n_3052), .CO(n_3093), .S(n_3092));
   HA_X1 i_2884 (.A(n_3038), .B(n_3031), .CO(n_3098), .S(n_3097));
   HA_X1 i_2888 (.A(n_3017), .B(n_3010), .CO(n_3103), .S(n_3102));
   HA_X1 i_2892 (.A(n_2938), .B(n_3084), .CO(n_3108), .S(n_3107));
   HA_X1 i_2896 (.A(n_3074), .B(n_2953), .CO(n_3113), .S(n_3112));
   HA_X1 i_2900 (.A(n_2943), .B(n_3089), .CO(n_3118), .S(n_3117));
   HA_X1 i_2904 (.A(n_2958), .B(n_3104), .CO(n_3123), .S(n_3122));
   HA_X1 i_2908 (.A(n_3094), .B(n_2968), .CO(n_3128), .S(n_3127));
   HA_X1 i_2912 (.A(n_3109), .B(n_2973), .CO(n_3133), .S(n_3132));
   HA_X1 i_2916 (.A(n_3119), .B(n_2983), .CO(n_3138), .S(n_3137));
   HA_X1 i_2920 (.A(n_3129), .B(n_2988), .CO(n_3143), .S(n_3142));
   HA_X1 i_2924 (.A(n_3139), .B(n_2993), .CO(n_3148), .S(n_3147));
   HA_X1 i_2928 (.A(n_2998), .B(n_3149), .CO(n_3153), .S(n_3152));
   HA_X1 i_2999 (.A(n_3060), .B(n_3053), .CO(n_3225), .S(n_3224));
   HA_X1 i_3003 (.A(n_3039), .B(n_3032), .CO(n_3230), .S(n_3229));
   HA_X1 i_3007 (.A(n_3018), .B(n_3011), .CO(n_3235), .S(n_3234));
   HA_X1 i_3011 (.A(n_3081), .B(n_3076), .CO(n_3240), .S(n_3239));
   HA_X1 i_3015 (.A(n_3219), .B(n_3212), .CO(n_3245), .S(n_3244));
   HA_X1 i_3019 (.A(n_3198), .B(n_3191), .CO(n_3250), .S(n_3249));
   HA_X1 i_3023 (.A(n_3177), .B(n_3170), .CO(n_3255), .S(n_3254));
   HA_X1 i_3027 (.A(n_3156), .B(n_3086), .CO(n_3260), .S(n_3259));
   HA_X1 i_3031 (.A(n_3231), .B(n_3226), .CO(n_3265), .S(n_3264));
   HA_X1 i_3035 (.A(n_3101), .B(n_3096), .CO(n_3270), .S(n_3269));
   HA_X1 i_3039 (.A(n_3241), .B(n_3116), .CO(n_3275), .S(n_3274));
   HA_X1 i_3043 (.A(n_3256), .B(n_3251), .CO(n_3280), .S(n_3279));
   HA_X1 i_3047 (.A(n_3261), .B(n_3121), .CO(n_3285), .S(n_3284));
   HA_X1 i_3051 (.A(n_3266), .B(n_3126), .CO(n_3290), .S(n_3289));
   HA_X1 i_3055 (.A(n_3131), .B(n_3136), .CO(n_3295), .S(n_3294));
   HA_X1 i_3059 (.A(n_3286), .B(n_3291), .CO(n_3300), .S(n_3299));
   HA_X1 i_3063 (.A(n_3146), .B(n_3296), .CO(n_3305), .S(n_3304));
   HA_X1 i_3067 (.A(n_3151), .B(n_3306), .CO(n_3310), .S(n_3309));
   HA_X1 i_3146 (.A(n_3206), .B(n_3199), .CO(n_3390), .S(n_3389));
   HA_X1 i_3150 (.A(n_3185), .B(n_3178), .CO(n_3395), .S(n_3394));
   HA_X1 i_3154 (.A(n_3164), .B(n_3157), .CO(n_3400), .S(n_3399));
   HA_X1 i_3158 (.A(n_3233), .B(n_3228), .CO(n_3405), .S(n_3404));
   HA_X1 i_3162 (.A(n_3369), .B(n_3362), .CO(n_3410), .S(n_3409));
   HA_X1 i_3166 (.A(n_3348), .B(n_3341), .CO(n_3415), .S(n_3414));
   HA_X1 i_3170 (.A(n_3327), .B(n_3320), .CO(n_3420), .S(n_3419));
   HA_X1 i_3174 (.A(n_3243), .B(n_3401), .CO(n_3425), .S(n_3424));
   HA_X1 i_3178 (.A(n_3391), .B(n_3383), .CO(n_3430), .S(n_3429));
   HA_X1 i_3182 (.A(n_3253), .B(n_3248), .CO(n_3435), .S(n_3434));
   HA_X1 i_3186 (.A(n_3273), .B(n_3268), .CO(n_3440), .S(n_3439));
   HA_X1 i_3190 (.A(n_3421), .B(n_3416), .CO(n_3445), .S(n_3444));
   HA_X1 i_3194 (.A(n_3278), .B(n_3436), .CO(n_3450), .S(n_3449));
   HA_X1 i_3198 (.A(n_3426), .B(n_3283), .CO(n_3455), .S(n_3454));
   HA_X1 i_3202 (.A(n_3288), .B(n_3446), .CO(n_3460), .S(n_3459));
   HA_X1 i_3206 (.A(n_3456), .B(n_3451), .CO(n_3465), .S(n_3464));
   HA_X1 i_3210 (.A(n_3303), .B(n_3461), .CO(n_3470), .S(n_3469));
   HA_X1 i_3214 (.A(n_3308), .B(n_3471), .CO(n_3475), .S(n_3474));
   HA_X1 i_3294 (.A(n_3370), .B(n_3363), .CO(n_3556), .S(n_3555));
   HA_X1 i_3298 (.A(n_3349), .B(n_3342), .CO(n_3561), .S(n_3560));
   HA_X1 i_3302 (.A(n_3328), .B(n_3321), .CO(n_3566), .S(n_3565));
   HA_X1 i_3306 (.A(n_3398), .B(n_3393), .CO(n_3571), .S(n_3570));
   HA_X1 i_3310 (.A(n_3549), .B(n_3542), .CO(n_3576), .S(n_3575));
   HA_X1 i_3314 (.A(n_3528), .B(n_3521), .CO(n_3581), .S(n_3580));
   HA_X1 i_3318 (.A(n_3507), .B(n_3500), .CO(n_3586), .S(n_3585));
   HA_X1 i_3322 (.A(n_3486), .B(n_3477), .CO(n_3591), .S(n_3590));
   HA_X1 i_3326 (.A(n_3567), .B(n_3562), .CO(n_3596), .S(n_3595));
   HA_X1 i_3330 (.A(n_3423), .B(n_3418), .CO(n_3601), .S(n_3600));
   HA_X1 i_3334 (.A(n_3408), .B(n_3572), .CO(n_3606), .S(n_3605));
   HA_X1 i_3338 (.A(n_3428), .B(n_3592), .CO(n_3611), .S(n_3610));
   HA_X1 i_3342 (.A(n_3582), .B(n_3577), .CO(n_3616), .S(n_3615));
   HA_X1 i_3346 (.A(n_3438), .B(n_3602), .CO(n_3621), .S(n_3620));
   HA_X1 i_3350 (.A(n_3448), .B(n_3607), .CO(n_3626), .S(n_3625));
   HA_X1 i_3354 (.A(n_3617), .B(n_3612), .CO(n_3631), .S(n_3630));
   HA_X1 i_3358 (.A(n_3622), .B(n_3463), .CO(n_3636), .S(n_3635));
   HA_X1 i_3362 (.A(n_3468), .B(n_3632), .CO(n_3641), .S(n_3640));
   HA_X1 i_3366 (.A(n_3473), .B(n_3642), .CO(n_3646), .S(n_3645));
   HA_X1 i_3442 (.A(n_3536), .B(n_3529), .CO(n_3723), .S(n_3722));
   HA_X1 i_3446 (.A(n_3515), .B(n_3508), .CO(n_3728), .S(n_3727));
   HA_X1 i_3450 (.A(n_3494), .B(n_3487), .CO(n_3733), .S(n_3732));
   HA_X1 i_3454 (.A(n_3569), .B(n_3564), .CO(n_3738), .S(n_3737));
   HA_X1 i_3458 (.A(n_3550), .B(n_3716), .CO(n_3743), .S(n_3742));
   HA_X1 i_3462 (.A(n_3702), .B(n_3695), .CO(n_3748), .S(n_3747));
   HA_X1 i_3466 (.A(n_3681), .B(n_3674), .CO(n_3753), .S(n_3752));
   HA_X1 i_3470 (.A(n_3660), .B(n_3653), .CO(n_3758), .S(n_3757));
   HA_X1 i_3474 (.A(n_3574), .B(n_3734), .CO(n_3763), .S(n_3762));
   HA_X1 i_3478 (.A(n_3724), .B(n_3589), .CO(n_3768), .S(n_3767));
   HA_X1 i_3482 (.A(n_3579), .B(n_3594), .CO(n_3773), .S(n_3772));
   HA_X1 i_3486 (.A(n_3604), .B(n_3599), .CO(n_3778), .S(n_3777));
   HA_X1 i_3490 (.A(n_3754), .B(n_3749), .CO(n_3783), .S(n_3782));
   HA_X1 i_3494 (.A(n_3609), .B(n_3769), .CO(n_3788), .S(n_3787));
   HA_X1 i_3498 (.A(n_3614), .B(n_3774), .CO(n_3793), .S(n_3792));
   HA_X1 i_3502 (.A(n_3779), .B(n_3624), .CO(n_3798), .S(n_3797));
   HA_X1 i_3506 (.A(n_3629), .B(n_3789), .CO(n_3803), .S(n_3802));
   HA_X1 i_3510 (.A(n_3634), .B(n_3799), .CO(n_3808), .S(n_3807));
   HA_X1 i_3514 (.A(n_3804), .B(n_3809), .CO(n_3813), .S(n_3812));
   HA_X1 i_3590 (.A(n_3710), .B(n_3703), .CO(n_3890), .S(n_3889));
   HA_X1 i_3594 (.A(n_3689), .B(n_3682), .CO(n_3895), .S(n_3894));
   HA_X1 i_3598 (.A(n_3668), .B(n_3661), .CO(n_3900), .S(n_3899));
   HA_X1 i_3602 (.A(n_3649), .B(n_3736), .CO(n_3905), .S(n_3904));
   HA_X1 i_3606 (.A(n_3726), .B(n_3717), .CO(n_3910), .S(n_3909));
   HA_X1 i_3610 (.A(n_3876), .B(n_3869), .CO(n_3915), .S(n_3914));
   HA_X1 i_3614 (.A(n_3855), .B(n_3848), .CO(n_3920), .S(n_3919));
   HA_X1 i_3618 (.A(n_3834), .B(n_3827), .CO(n_3925), .S(n_3924));
   HA_X1 i_3622 (.A(n_3741), .B(n_3901), .CO(n_3930), .S(n_3929));
   HA_X1 i_3626 (.A(n_3891), .B(n_3761), .CO(n_3935), .S(n_3934));
   HA_X1 i_3630 (.A(n_3751), .B(n_3746), .CO(n_3940), .S(n_3939));
   HA_X1 i_3634 (.A(n_3906), .B(n_3771), .CO(n_3945), .S(n_3944));
   HA_X1 i_3638 (.A(n_3926), .B(n_3921), .CO(n_3950), .S(n_3949));
   HA_X1 i_3642 (.A(n_3776), .B(n_3941), .CO(n_3955), .S(n_3954));
   HA_X1 i_3646 (.A(n_3931), .B(n_3786), .CO(n_3960), .S(n_3959));
   HA_X1 i_3650 (.A(n_3946), .B(n_3791), .CO(n_3965), .S(n_3964));
   HA_X1 i_3654 (.A(n_3951), .B(n_3961), .CO(n_3970), .S(n_3969));
   HA_X1 i_3658 (.A(n_3801), .B(n_3966), .CO(n_3975), .S(n_3974));
   HA_X1 i_3662 (.A(n_3971), .B(n_3811), .CO(n_3980), .S(n_3979));
   HA_X1 i_3738 (.A(n_3877), .B(n_3870), .CO(n_4057), .S(n_4056));
   HA_X1 i_3742 (.A(n_3856), .B(n_3849), .CO(n_4062), .S(n_4061));
   HA_X1 i_3746 (.A(n_3835), .B(n_3828), .CO(n_4067), .S(n_4066));
   HA_X1 i_3750 (.A(n_3903), .B(n_3898), .CO(n_4072), .S(n_4071));
   HA_X1 i_3754 (.A(n_4050), .B(n_4043), .CO(n_4077), .S(n_4076));
   HA_X1 i_3758 (.A(n_4029), .B(n_4022), .CO(n_4082), .S(n_4081));
   HA_X1 i_3762 (.A(n_4008), .B(n_4001), .CO(n_4087), .S(n_4086));
   HA_X1 i_3766 (.A(n_3985), .B(n_3908), .CO(n_4092), .S(n_4091));
   HA_X1 i_3770 (.A(n_4063), .B(n_4058), .CO(n_4097), .S(n_4096));
   HA_X1 i_3774 (.A(n_3923), .B(n_3918), .CO(n_4102), .S(n_4101));
   HA_X1 i_3778 (.A(n_4073), .B(n_3938), .CO(n_4107), .S(n_4106));
   HA_X1 i_3782 (.A(n_4088), .B(n_4083), .CO(n_4112), .S(n_4111));
   HA_X1 i_3786 (.A(n_4093), .B(n_3948), .CO(n_4117), .S(n_4116));
   HA_X1 i_3790 (.A(n_4103), .B(n_4098), .CO(n_4122), .S(n_4121));
   HA_X1 i_3794 (.A(n_4108), .B(n_3963), .CO(n_4127), .S(n_4126));
   HA_X1 i_3798 (.A(n_4113), .B(n_4118), .CO(n_4132), .S(n_4131));
   HA_X1 i_3802 (.A(n_4123), .B(n_4128), .CO(n_4137), .S(n_4136));
   HA_X1 i_3806 (.A(n_4133), .B(n_3978), .CO(n_4142), .S(n_4141));
   HA_X1 i_3874 (.A(n_384), .B(n_4044), .CO(n_4211), .S(n_4210));
   HA_X1 i_3878 (.A(n_4030), .B(n_4023), .CO(n_4216), .S(n_4215));
   HA_X1 i_3882 (.A(n_4009), .B(n_4002), .CO(n_4221), .S(n_4220));
   HA_X1 i_3886 (.A(n_3986), .B(n_4070), .CO(n_4226), .S(n_4225));
   HA_X1 i_3890 (.A(n_4060), .B(n_4051), .CO(n_4231), .S(n_4230));
   HA_X1 i_3894 (.A(n_4198), .B(n_4191), .CO(n_4236), .S(n_4235));
   HA_X1 i_3898 (.A(n_4177), .B(n_4170), .CO(n_4241), .S(n_4240));
   HA_X1 i_3902 (.A(n_4156), .B(n_4147), .CO(n_4246), .S(n_4245));
   HA_X1 i_3906 (.A(n_4222), .B(n_4217), .CO(n_4251), .S(n_4250));
   HA_X1 i_3910 (.A(n_4090), .B(n_4085), .CO(n_4256), .S(n_4255));
   HA_X1 i_3914 (.A(n_4232), .B(n_4227), .CO(n_4261), .S(n_4260));
   HA_X1 i_3918 (.A(n_4100), .B(n_4095), .CO(n_4266), .S(n_4265));
   HA_X1 i_3922 (.A(n_4242), .B(n_4237), .CO(n_4271), .S(n_4270));
   HA_X1 i_3926 (.A(n_4257), .B(n_4252), .CO(n_4276), .S(n_4275));
   HA_X1 i_3930 (.A(n_4120), .B(n_4267), .CO(n_4281), .S(n_4280));
   HA_X1 i_3934 (.A(n_4125), .B(n_4272), .CO(n_4286), .S(n_4285));
   HA_X1 i_3938 (.A(n_4277), .B(n_4135), .CO(n_4291), .S(n_4290));
   HA_X1 i_3942 (.A(n_4287), .B(n_4140), .CO(n_4296), .S(n_4295));
   HA_X1 i_4011 (.A(n_4206), .B(n_4199), .CO(n_4366), .S(n_4365));
   HA_X1 i_4015 (.A(n_4185), .B(n_4178), .CO(n_4371), .S(n_4370));
   HA_X1 i_4019 (.A(n_4164), .B(n_4157), .CO(n_4376), .S(n_4375));
   HA_X1 i_4023 (.A(n_4224), .B(n_4219), .CO(n_4381), .S(n_4380));
   HA_X1 i_4027 (.A(n_4358), .B(n_4352), .CO(n_4386), .S(n_4385));
   HA_X1 i_4031 (.A(n_4338), .B(n_4331), .CO(n_4391), .S(n_4390));
   HA_X1 i_4035 (.A(n_4317), .B(n_4310), .CO(n_4396), .S(n_4395));
   HA_X1 i_4039 (.A(n_4229), .B(n_4377), .CO(n_4401), .S(n_4400));
   HA_X1 i_4043 (.A(n_4367), .B(n_4244), .CO(n_4406), .S(n_4405));
   HA_X1 i_4047 (.A(n_4234), .B(n_4249), .CO(n_4411), .S(n_4410));
   HA_X1 i_4051 (.A(n_4259), .B(n_4254), .CO(n_4416), .S(n_4415));
   HA_X1 i_4055 (.A(n_4392), .B(n_4387), .CO(n_4421), .S(n_4420));
   HA_X1 i_4059 (.A(n_4407), .B(n_4402), .CO(n_4426), .S(n_4425));
   HA_X1 i_4063 (.A(n_4412), .B(n_4274), .CO(n_4431), .S(n_4430));
   HA_X1 i_4067 (.A(n_4279), .B(n_4422), .CO(n_4436), .S(n_4435));
   HA_X1 i_4071 (.A(n_4427), .B(n_4432), .CO(n_4441), .S(n_4440));
   HA_X1 i_4075 (.A(n_4437), .B(n_4294), .CO(n_4446), .S(n_4445));
   HA_X1 i_4144 (.A(n_4353), .B(n_4346), .CO(n_4516), .S(n_4515));
   HA_X1 i_4148 (.A(n_4332), .B(n_4325), .CO(n_4521), .S(n_4520));
   HA_X1 i_4152 (.A(n_4311), .B(n_4302), .CO(n_4526), .S(n_4525));
   HA_X1 i_4156 (.A(n_4374), .B(n_4369), .CO(n_4531), .S(n_4530));
   HA_X1 i_4160 (.A(n_4502), .B(n_4495), .CO(n_4536), .S(n_4535));
   HA_X1 i_4164 (.A(n_4481), .B(n_4474), .CO(n_4541), .S(n_4540));
   HA_X1 i_4168 (.A(n_4460), .B(n_4451), .CO(n_4546), .S(n_4545));
   HA_X1 i_4172 (.A(n_4527), .B(n_4522), .CO(n_4551), .S(n_4550));
   HA_X1 i_4176 (.A(n_4399), .B(n_4394), .CO(n_4556), .S(n_4555));
   HA_X1 i_4180 (.A(n_4532), .B(n_4409), .CO(n_4561), .S(n_4560));
   HA_X1 i_4184 (.A(n_4547), .B(n_4542), .CO(n_4566), .S(n_4565));
   HA_X1 i_4188 (.A(n_4414), .B(n_4557), .CO(n_4571), .S(n_4570));
   HA_X1 i_4192 (.A(n_4419), .B(n_4424), .CO(n_4576), .S(n_4575));
   HA_X1 i_4196 (.A(n_4429), .B(n_4567), .CO(n_4581), .S(n_4580));
   HA_X1 i_4200 (.A(n_4572), .B(n_4577), .CO(n_4586), .S(n_4585));
   HA_X1 i_4204 (.A(n_4444), .B(n_4582), .CO(n_4591), .S(n_4590));
   HA_X1 i_4265 (.A(n_383), .B(n_4503), .CO(n_4653), .S(n_4652));
   HA_X1 i_4269 (.A(n_4489), .B(n_4482), .CO(n_4658), .S(n_4657));
   HA_X1 i_4273 (.A(n_4468), .B(n_4461), .CO(n_4663), .S(n_4662));
   HA_X1 i_4277 (.A(n_4524), .B(n_4519), .CO(n_4668), .S(n_4667));
   HA_X1 i_4281 (.A(n_4647), .B(n_4640), .CO(n_4673), .S(n_4672));
   HA_X1 i_4285 (.A(n_4626), .B(n_4619), .CO(n_4678), .S(n_4677));
   HA_X1 i_4289 (.A(n_4605), .B(n_4596), .CO(n_4683), .S(n_4682));
   HA_X1 i_4293 (.A(n_4664), .B(n_4659), .CO(n_4688), .S(n_4687));
   HA_X1 i_4297 (.A(n_4544), .B(n_4539), .CO(n_4693), .S(n_4692));
   HA_X1 i_4301 (.A(n_4549), .B(n_4669), .CO(n_4698), .S(n_4697));
   HA_X1 i_4305 (.A(n_4554), .B(n_4684), .CO(n_4703), .S(n_4702));
   HA_X1 i_4309 (.A(n_4674), .B(n_4564), .CO(n_4708), .S(n_4707));
   HA_X1 i_4313 (.A(n_4689), .B(n_4569), .CO(n_4713), .S(n_4712));
   HA_X1 i_4317 (.A(n_4574), .B(n_4704), .CO(n_4718), .S(n_4717));
   HA_X1 i_4321 (.A(n_4579), .B(n_4714), .CO(n_4723), .S(n_4722));
   HA_X1 i_4325 (.A(n_4589), .B(n_4719), .CO(n_4728), .S(n_4727));
   HA_X1 i_4387 (.A(n_4648), .B(n_4641), .CO(n_4791), .S(n_4790));
   HA_X1 i_4391 (.A(n_4627), .B(n_4620), .CO(n_4796), .S(n_4795));
   HA_X1 i_4395 (.A(n_4606), .B(n_4597), .CO(n_4801), .S(n_4800));
   HA_X1 i_4399 (.A(n_4661), .B(n_4656), .CO(n_4806), .S(n_4805));
   HA_X1 i_4403 (.A(n_4777), .B(n_4770), .CO(n_4811), .S(n_4810));
   HA_X1 i_4407 (.A(n_4756), .B(n_4749), .CO(n_4816), .S(n_4815));
   HA_X1 i_4411 (.A(n_4733), .B(n_4671), .CO(n_4821), .S(n_4820));
   HA_X1 i_4415 (.A(n_4797), .B(n_4792), .CO(n_4826), .S(n_4825));
   HA_X1 i_4419 (.A(n_4676), .B(n_4686), .CO(n_4831), .S(n_4830));
   HA_X1 i_4423 (.A(n_4696), .B(n_4691), .CO(n_4836), .S(n_4835));
   HA_X1 i_4427 (.A(n_4812), .B(n_4822), .CO(n_4841), .S(n_4840));
   HA_X1 i_4431 (.A(n_4827), .B(n_4706), .CO(n_4846), .S(n_4845));
   HA_X1 i_4435 (.A(n_4837), .B(n_4711), .CO(n_4851), .S(n_4850));
   HA_X1 i_4439 (.A(n_4716), .B(n_4847), .CO(n_4856), .S(n_4855));
   HA_X1 i_4443 (.A(n_4852), .B(n_4726), .CO(n_4861), .S(n_4860));
   HA_X1 i_4505 (.A(n_4778), .B(n_4771), .CO(n_4924), .S(n_4923));
   HA_X1 i_4509 (.A(n_4757), .B(n_4750), .CO(n_4929), .S(n_4928));
   HA_X1 i_4513 (.A(n_4734), .B(n_4799), .CO(n_4934), .S(n_4933));
   HA_X1 i_4517 (.A(n_4917), .B(n_4910), .CO(n_4939), .S(n_4938));
   HA_X1 i_4521 (.A(n_4896), .B(n_4889), .CO(n_4944), .S(n_4943));
   HA_X1 i_4525 (.A(n_4875), .B(n_4866), .CO(n_4949), .S(n_4948));
   HA_X1 i_4529 (.A(n_4930), .B(n_4925), .CO(n_4954), .S(n_4953));
   HA_X1 i_4533 (.A(n_4814), .B(n_4809), .CO(n_4959), .S(n_4958));
   HA_X1 i_4537 (.A(n_4829), .B(n_4824), .CO(n_4964), .S(n_4963));
   HA_X1 i_4541 (.A(n_4945), .B(n_4940), .CO(n_4969), .S(n_4968));
   HA_X1 i_4545 (.A(n_4960), .B(n_4955), .CO(n_4974), .S(n_4973));
   HA_X1 i_4549 (.A(n_4844), .B(n_4965), .CO(n_4979), .S(n_4978));
   HA_X1 i_4553 (.A(n_4970), .B(n_4975), .CO(n_4984), .S(n_4983));
   HA_X1 i_4557 (.A(n_4980), .B(n_4859), .CO(n_4989), .S(n_4988));
   HA_X1 i_4611 (.A(n_382), .B(n_4911), .CO(n_5044), .S(n_5043));
   HA_X1 i_4615 (.A(n_4897), .B(n_4890), .CO(n_5049), .S(n_5048));
   HA_X1 i_4619 (.A(n_4876), .B(n_4867), .CO(n_5054), .S(n_5053));
   HA_X1 i_4623 (.A(n_4927), .B(n_4918), .CO(n_5059), .S(n_5058));
   HA_X1 i_4627 (.A(n_5031), .B(n_5024), .CO(n_5064), .S(n_5063));
   HA_X1 i_4631 (.A(n_5010), .B(n_5003), .CO(n_5069), .S(n_5068));
   HA_X1 i_4635 (.A(n_4937), .B(n_5055), .CO(n_5074), .S(n_5073));
   HA_X1 i_4639 (.A(n_5045), .B(n_4947), .CO(n_5079), .S(n_5078));
   HA_X1 i_4643 (.A(n_4952), .B(n_5060), .CO(n_5084), .S(n_5083));
   HA_X1 i_4647 (.A(n_5070), .B(n_5065), .CO(n_5089), .S(n_5088));
   HA_X1 i_4651 (.A(n_5080), .B(n_5075), .CO(n_5094), .S(n_5093));
   HA_X1 i_4655 (.A(n_4972), .B(n_5085), .CO(n_5099), .S(n_5098));
   HA_X1 i_4659 (.A(n_5090), .B(n_4982), .CO(n_5104), .S(n_5103));
   HA_X1 i_4663 (.A(n_5100), .B(n_4987), .CO(n_5109), .S(n_5108));
   HA_X1 i_4718 (.A(n_5039), .B(n_5032), .CO(n_5165), .S(n_5164));
   HA_X1 i_4722 (.A(n_5018), .B(n_5011), .CO(n_5170), .S(n_5169));
   HA_X1 i_4726 (.A(n_4995), .B(n_5052), .CO(n_5175), .S(n_5174));
   HA_X1 i_4730 (.A(n_5157), .B(n_5151), .CO(n_5180), .S(n_5179));
   HA_X1 i_4734 (.A(n_5137), .B(n_5130), .CO(n_5185), .S(n_5184));
   HA_X1 i_4738 (.A(n_5114), .B(n_5057), .CO(n_5190), .S(n_5189));
   HA_X1 i_4742 (.A(n_5166), .B(n_5072), .CO(n_5195), .S(n_5194));
   HA_X1 i_4746 (.A(n_5062), .B(n_5176), .CO(n_5200), .S(n_5199));
   HA_X1 i_4750 (.A(n_5077), .B(n_5186), .CO(n_5205), .S(n_5204));
   HA_X1 i_4754 (.A(n_5191), .B(n_5087), .CO(n_5210), .S(n_5209));
   HA_X1 i_4758 (.A(n_5092), .B(n_5201), .CO(n_5215), .S(n_5214));
   HA_X1 i_4762 (.A(n_5206), .B(n_5211), .CO(n_5220), .S(n_5219));
   HA_X1 i_4766 (.A(n_5216), .B(n_5107), .CO(n_5225), .S(n_5224));
   HA_X1 i_4821 (.A(n_5152), .B(n_5145), .CO(n_5281), .S(n_5280));
   HA_X1 i_4825 (.A(n_5131), .B(n_5124), .CO(n_5286), .S(n_5285));
   HA_X1 i_4829 (.A(n_5173), .B(n_5168), .CO(n_5291), .S(n_5290));
   HA_X1 i_4833 (.A(n_5267), .B(n_5260), .CO(n_5296), .S(n_5295));
   HA_X1 i_4837 (.A(n_5246), .B(n_5239), .CO(n_5301), .S(n_5300));
   HA_X1 i_4841 (.A(n_5178), .B(n_5287), .CO(n_5306), .S(n_5305));
   HA_X1 i_4845 (.A(n_5188), .B(n_5183), .CO(n_5311), .S(n_5310));
   HA_X1 i_4849 (.A(n_5198), .B(n_5193), .CO(n_5316), .S(n_5315));
   HA_X1 i_4853 (.A(n_5297), .B(n_5203), .CO(n_5321), .S(n_5320));
   HA_X1 i_4857 (.A(n_5307), .B(n_5208), .CO(n_5326), .S(n_5325));
   HA_X1 i_4861 (.A(n_5213), .B(n_5322), .CO(n_5331), .S(n_5330));
   HA_X1 i_4865 (.A(n_5327), .B(n_5223), .CO(n_5336), .S(n_5335));
   HA_X1 i_4912 (.A(n_447), .B(n_5268), .CO(n_5384), .S(n_5383));
   HA_X1 i_4916 (.A(n_5254), .B(n_5247), .CO(n_5389), .S(n_5388));
   HA_X1 i_4920 (.A(n_5231), .B(n_5289), .CO(n_5394), .S(n_5393));
   HA_X1 i_4924 (.A(n_5275), .B(n_5378), .CO(n_5399), .S(n_5398));
   HA_X1 i_4928 (.A(n_5364), .B(n_5357), .CO(n_5404), .S(n_5403));
   HA_X1 i_4932 (.A(n_5341), .B(n_5390), .CO(n_5409), .S(n_5408));
   HA_X1 i_4936 (.A(n_5304), .B(n_5299), .CO(n_5414), .S(n_5413));
   HA_X1 i_4940 (.A(n_5395), .B(n_5309), .CO(n_5419), .S(n_5418));
   HA_X1 i_4944 (.A(n_5400), .B(n_5314), .CO(n_5424), .S(n_5423));
   HA_X1 i_4948 (.A(n_5410), .B(n_5319), .CO(n_5429), .S(n_5428));
   HA_X1 i_4952 (.A(n_5324), .B(n_5425), .CO(n_5434), .S(n_5433));
   HA_X1 i_4956 (.A(n_5430), .B(n_5334), .CO(n_5439), .S(n_5438));
   HA_X1 i_5004 (.A(n_5379), .B(n_5372), .CO(n_5488), .S(n_5487));
   HA_X1 i_5008 (.A(n_5358), .B(n_5351), .CO(n_5493), .S(n_5492));
   HA_X1 i_5012 (.A(n_5392), .B(n_5387), .CO(n_5498), .S(n_5497));
   HA_X1 i_5016 (.A(n_5474), .B(n_5467), .CO(n_5503), .S(n_5502));
   HA_X1 i_5020 (.A(n_5453), .B(n_5444), .CO(n_5508), .S(n_5507));
   HA_X1 i_5024 (.A(n_5494), .B(n_5489), .CO(n_5513), .S(n_5512));
   HA_X1 i_5028 (.A(n_5402), .B(n_5499), .CO(n_5518), .S(n_5517));
   HA_X1 i_5032 (.A(n_5412), .B(n_5509), .CO(n_5523), .S(n_5522));
   HA_X1 i_5036 (.A(n_5514), .B(n_5422), .CO(n_5528), .S(n_5527));
   HA_X1 i_5040 (.A(n_5427), .B(n_5524), .CO(n_5533), .S(n_5532));
   HA_X1 i_5044 (.A(n_5529), .B(n_5437), .CO(n_5538), .S(n_5537));
   HA_X1 i_5092 (.A(n_5475), .B(n_5468), .CO(n_5587), .S(n_5586));
   HA_X1 i_5096 (.A(n_5454), .B(n_5445), .CO(n_5592), .S(n_5591));
   HA_X1 i_5100 (.A(n_5491), .B(n_5580), .CO(n_5597), .S(n_5596));
   HA_X1 i_5104 (.A(n_5566), .B(n_5559), .CO(n_5602), .S(n_5601));
   HA_X1 i_5108 (.A(n_5543), .B(n_5593), .CO(n_5607), .S(n_5606));
   HA_X1 i_5112 (.A(n_5506), .B(n_5501), .CO(n_5612), .S(n_5611));
   HA_X1 i_5116 (.A(n_5516), .B(n_5603), .CO(n_5617), .S(n_5616));
   HA_X1 i_5120 (.A(n_5521), .B(n_5613), .CO(n_5622), .S(n_5621));
   HA_X1 i_5124 (.A(n_5526), .B(n_5618), .CO(n_5627), .S(n_5626));
   HA_X1 i_5128 (.A(n_5623), .B(n_5536), .CO(n_5632), .S(n_5631));
   HA_X1 i_5168 (.A(n_543), .B(n_5574), .CO(n_5673), .S(n_5672));
   HA_X1 i_5172 (.A(n_5560), .B(n_5553), .CO(n_5678), .S(n_5677));
   HA_X1 i_5176 (.A(n_5590), .B(n_5581), .CO(n_5683), .S(n_5682));
   HA_X1 i_5180 (.A(n_5660), .B(n_5653), .CO(n_5688), .S(n_5687));
   HA_X1 i_5184 (.A(n_5637), .B(n_5595), .CO(n_5693), .S(n_5692));
   HA_X1 i_5188 (.A(n_5674), .B(n_5605), .CO(n_5698), .S(n_5697));
   HA_X1 i_5192 (.A(n_5684), .B(n_5610), .CO(n_5703), .S(n_5702));
   HA_X1 i_5196 (.A(n_5689), .B(n_5694), .CO(n_5708), .S(n_5707));
   HA_X1 i_5200 (.A(n_5620), .B(n_5704), .CO(n_5713), .S(n_5712));
   HA_X1 i_5204 (.A(n_5709), .B(n_5630), .CO(n_5718), .S(n_5717));
   HA_X1 i_5245 (.A(n_5668), .B(n_5661), .CO(n_5760), .S(n_5759));
   HA_X1 i_5249 (.A(n_5647), .B(n_5638), .CO(n_5765), .S(n_5764));
   HA_X1 i_5253 (.A(n_5676), .B(n_5752), .CO(n_1), .S(n_0));
   HA_X1 i_5257 (.A(n_5739), .B(n_5732), .CO(n_3), .S(n_2));
   HA_X1 i_5261 (.A(n_5766), .B(n_5761), .CO(n_5), .S(n_4));
   HA_X1 i_5265 (.A(n_5686), .B(n_5701), .CO(n_7), .S(n_6));
   HA_X1 i_5269 (.A(n_381), .B(n_380), .CO(n_9), .S(n_8));
   HA_X1 i_5273 (.A(n_379), .B(n_378), .CO(n_11), .S(n_10));
   HA_X1 i_5277 (.A(n_377), .B(n_5716), .CO(n_13), .S(n_12));
   HA_X1 i_5318 (.A(n_5747), .B(n_5740), .CO(n_15), .S(n_14));
   HA_X1 i_5322 (.A(n_5724), .B(n_5763), .CO(n_17), .S(n_16));
   HA_X1 i_5326 (.A(n_376), .B(n_375), .CO(n_19), .S(n_18));
   HA_X1 i_5330 (.A(n_374), .B(n_373), .CO(n_21), .S(n_20));
   HA_X1 i_5334 (.A(n_372), .B(n_371), .CO(n_23), .S(n_22));
   HA_X1 i_5338 (.A(n_370), .B(n_369), .CO(n_25), .S(n_24));
   HA_X1 i_5342 (.A(n_368), .B(n_367), .CO(n_27), .S(n_26));
   HA_X1 i_5346 (.A(n_366), .B(n_365), .CO(n_29), .S(n_28));
   HA_X1 i_5379 (.A(n_639), .B(n_364), .CO(n_31), .S(n_30));
   HA_X1 i_5383 (.A(n_363), .B(n_362), .CO(n_33), .S(n_32));
   HA_X1 i_5387 (.A(n_361), .B(n_360), .CO(n_35), .S(n_34));
   HA_X1 i_5391 (.A(n_359), .B(n_358), .CO(n_37), .S(n_36));
   HA_X1 i_5395 (.A(n_357), .B(n_356), .CO(n_39), .S(n_38));
   HA_X1 i_5399 (.A(n_355), .B(n_354), .CO(n_41), .S(n_40));
   HA_X1 i_5403 (.A(n_353), .B(n_352), .CO(n_43), .S(n_42));
   HA_X1 i_5407 (.A(n_351), .B(n_350), .CO(n_45), .S(n_44));
   HA_X1 i_5441 (.A(n_349), .B(n_348), .CO(n_47), .S(n_46));
   HA_X1 i_5445 (.A(n_347), .B(n_346), .CO(n_49), .S(n_48));
   HA_X1 i_5449 (.A(n_345), .B(n_344), .CO(n_51), .S(n_50));
   HA_X1 i_5453 (.A(n_343), .B(n_342), .CO(n_53), .S(n_52));
   HA_X1 i_5457 (.A(n_341), .B(n_340), .CO(n_55), .S(n_54));
   HA_X1 i_5461 (.A(n_339), .B(n_338), .CO(n_57), .S(n_56));
   HA_X1 i_5465 (.A(n_337), .B(n_336), .CO(n_59), .S(n_58));
   HA_X1 i_5499 (.A(n_335), .B(n_334), .CO(n_61), .S(n_60));
   HA_X1 i_5503 (.A(n_333), .B(n_332), .CO(n_63), .S(n_62));
   HA_X1 i_5507 (.A(n_331), .B(n_330), .CO(n_65), .S(n_64));
   HA_X1 i_5511 (.A(n_329), .B(n_328), .CO(n_67), .S(n_66));
   HA_X1 i_5515 (.A(n_327), .B(n_326), .CO(n_69), .S(n_68));
   HA_X1 i_5519 (.A(n_325), .B(n_324), .CO(n_71), .S(n_70));
   HA_X1 i_5545 (.A(n_735), .B(n_323), .CO(n_73), .S(n_72));
   HA_X1 i_5549 (.A(n_322), .B(n_321), .CO(n_75), .S(n_74));
   HA_X1 i_5553 (.A(n_320), .B(n_319), .CO(n_77), .S(n_76));
   HA_X1 i_5557 (.A(n_318), .B(n_317), .CO(n_79), .S(n_78));
   HA_X1 i_5561 (.A(n_316), .B(n_315), .CO(n_81), .S(n_80));
   HA_X1 i_5565 (.A(n_314), .B(n_313), .CO(n_83), .S(n_82));
   HA_X1 i_5592 (.A(n_312), .B(n_311), .CO(n_85), .S(n_84));
   HA_X1 i_5596 (.A(n_310), .B(n_309), .CO(n_87), .S(n_86));
   HA_X1 i_5600 (.A(n_308), .B(n_307), .CO(n_89), .S(n_88));
   HA_X1 i_5604 (.A(n_306), .B(n_305), .CO(n_91), .S(n_90));
   HA_X1 i_5608 (.A(n_304), .B(n_303), .CO(n_93), .S(n_92));
   HA_X1 i_5635 (.A(n_302), .B(n_301), .CO(n_95), .S(n_94));
   HA_X1 i_5639 (.A(n_300), .B(n_299), .CO(n_97), .S(n_96));
   HA_X1 i_5643 (.A(n_298), .B(n_297), .CO(n_99), .S(n_98));
   HA_X1 i_5647 (.A(n_296), .B(n_295), .CO(n_101), .S(n_100));
   HA_X1 i_5666 (.A(n_831), .B(n_294), .CO(n_103), .S(n_102));
   HA_X1 i_5670 (.A(n_293), .B(n_292), .CO(n_105), .S(n_104));
   HA_X1 i_5674 (.A(n_291), .B(n_290), .CO(n_107), .S(n_106));
   HA_X1 i_5678 (.A(n_289), .B(n_288), .CO(n_109), .S(n_108));
   HA_X1 i_5698 (.A(n_287), .B(n_286), .CO(n_111), .S(n_110));
   HA_X1 i_5702 (.A(n_285), .B(n_284), .CO(n_113), .S(n_112));
   HA_X1 i_5706 (.A(n_283), .B(n_282), .CO(n_115), .S(n_114));
   HA_X1 i_5726 (.A(n_281), .B(n_280), .CO(n_117), .S(n_116));
   HA_X1 i_5730 (.A(n_279), .B(n_278), .CO(n_119), .S(n_118));
   HA_X1 i_5742 (.A(n_927), .B(n_277), .CO(n_121), .S(n_120));
   HA_X1 i_5746 (.A(n_276), .B(n_275), .CO(n_123), .S(n_122));
   HA_X1 i_5758 (.A(n_274), .B(n_273), .CO(n_125), .S(n_124));
   HA_X1 i_5762 (.A(n_1022), .B(n_991), .CO(n_127), .S(n_126));
   HA_X1 i_5778 (.A(n_1034), .B(n_1029), .CO(n_129), .S(n_128));
   HA_X1 i_5782 (.A(n_1039), .B(n_1052), .CO(n_131), .S(n_130));
   HA_X1 i_5786 (.A(n_1073), .B(n_1070), .CO(n_133), .S(n_132));
   HA_X1 i_5790 (.A(n_1102), .B(n_1099), .CO(n_135), .S(n_134));
   HA_X1 i_5794 (.A(n_1133), .B(n_1136), .CO(n_137), .S(n_136));
   HA_X1 i_5798 (.A(n_1171), .B(n_1174), .CO(n_139), .S(n_138));
   HA_X1 i_5802 (.A(n_1220), .B(n_1217), .CO(n_141), .S(n_140));
   HA_X1 i_5806 (.A(n_1271), .B(n_1268), .CO(n_143), .S(n_142));
   HA_X1 i_5810 (.A(n_1323), .B(n_1326), .CO(n_145), .S(n_144));
   HA_X1 i_5814 (.A(n_1386), .B(n_1389), .CO(n_147), .S(n_146));
   HA_X1 i_5818 (.A(n_1454), .B(n_1457), .CO(n_149), .S(n_148));
   HA_X1 i_5822 (.A(n_1526), .B(n_1529), .CO(n_151), .S(n_150));
   HA_X1 i_5826 (.A(n_1606), .B(n_1609), .CO(n_153), .S(n_152));
   HA_X1 i_5830 (.A(n_1691), .B(n_1694), .CO(n_155), .S(n_154));
   HA_X1 i_5834 (.A(n_1780), .B(n_1783), .CO(n_157), .S(n_156));
   HA_X1 i_5838 (.A(n_1784), .B(n_1880), .CO(n_159), .S(n_158));
   HA_X1 i_5842 (.A(n_1881), .B(n_1982), .CO(n_161), .S(n_160));
   HA_X1 i_5846 (.A(n_2085), .B(n_2088), .CO(n_163), .S(n_162));
   HA_X1 i_5850 (.A(n_2089), .B(n_2202), .CO(n_165), .S(n_164));
   HA_X1 i_5854 (.A(n_2203), .B(n_2321), .CO(n_167), .S(n_166));
   HA_X1 i_5858 (.A(n_2322), .B(n_2444), .CO(n_169), .S(n_168));
   HA_X1 i_5862 (.A(n_2445), .B(n_2575), .CO(n_171), .S(n_170));
   HA_X1 i_5866 (.A(n_2708), .B(n_2711), .CO(n_173), .S(n_172));
   HA_X1 i_5870 (.A(n_2712), .B(n_2851), .CO(n_175), .S(n_174));
   HA_X1 i_5874 (.A(n_2852), .B(n_2999), .CO(n_177), .S(n_176));
   HA_X1 i_5878 (.A(n_3000), .B(n_3152), .CO(n_179), .S(n_178));
   HA_X1 i_5882 (.A(n_3153), .B(n_3309), .CO(n_181), .S(n_180));
   HA_X1 i_5886 (.A(n_3310), .B(n_3474), .CO(n_183), .S(n_182));
   HA_X1 i_5890 (.A(n_3475), .B(n_3645), .CO(n_185), .S(n_184));
   HA_X1 i_5894 (.A(n_3646), .B(n_3814), .CO(n_187), .S(n_186));
   HA_X1 i_5898 (.A(n_3816), .B(n_3981), .CO(n_189), .S(n_188));
   HA_X1 i_5902 (.A(n_3983), .B(n_4143), .CO(n_191), .S(n_190));
   HA_X1 i_5906 (.A(n_4297), .B(n_4145), .CO(n_193), .S(n_192));
   HA_X1 i_5910 (.A(n_4299), .B(n_4447), .CO(n_195), .S(n_194));
   HA_X1 i_5914 (.A(n_4449), .B(n_4592), .CO(n_197), .S(n_196));
   HA_X1 i_5918 (.A(n_4594), .B(n_4729), .CO(n_199), .S(n_198));
   HA_X1 i_5922 (.A(n_4731), .B(n_4862), .CO(n_201), .S(n_200));
   HA_X1 i_5926 (.A(n_4864), .B(n_4990), .CO(n_203), .S(n_202));
   HA_X1 i_5930 (.A(n_4992), .B(n_5110), .CO(n_205), .S(n_204));
   HA_X1 i_5934 (.A(n_5112), .B(n_5226), .CO(n_207), .S(n_206));
   HA_X1 i_5938 (.A(n_5228), .B(n_5337), .CO(n_209), .S(n_208));
   HA_X1 i_5942 (.A(n_5339), .B(n_5440), .CO(n_211), .S(n_210));
   HA_X1 i_5946 (.A(n_5442), .B(n_5539), .CO(n_213), .S(n_212));
   HA_X1 i_5950 (.A(n_5541), .B(n_5633), .CO(n_215), .S(n_214));
   HA_X1 i_5954 (.A(n_5635), .B(n_5719), .CO(n_217), .S(n_216));
   HA_X1 i_5958 (.A(n_5721), .B(n_272), .CO(n_219), .S(n_218));
   HA_X1 i_5962 (.A(n_271), .B(n_270), .CO(n_221), .S(n_220));
   HA_X1 i_5966 (.A(n_269), .B(n_268), .CO(n_223), .S(n_222));
   HA_X1 i_5970 (.A(n_267), .B(n_266), .CO(n_225), .S(n_224));
   HA_X1 i_5974 (.A(n_265), .B(n_264), .CO(n_227), .S(n_226));
   HA_X1 i_5978 (.A(n_263), .B(n_262), .CO(n_229), .S(n_228));
   HA_X1 i_5982 (.A(n_261), .B(n_260), .CO(n_231), .S(n_230));
   HA_X1 i_5986 (.A(n_259), .B(n_258), .CO(n_233), .S(n_232));
   HA_X1 i_5990 (.A(n_257), .B(n_256), .CO(n_235), .S(n_234));
   HA_X1 i_5994 (.A(n_255), .B(n_254), .CO(n_237), .S(n_236));
   HA_X1 i_5998 (.A(n_253), .B(n_252), .CO(n_239), .S(n_238));
   HA_X1 i_6002 (.A(n_251), .B(n_250), .CO(n_241), .S(n_240));
   HA_X1 i_6006 (.A(n_249), .B(n_248), .CO(n_243), .S(n_242));
   HA_X1 i_6010 (.A(n_247), .B(n_246), .CO(n_245), .S(n_244));
   INV_X1 i_0 (.A(n_385), .ZN(n_246));
   AOI21_X1 i_1 (.A(n_125), .B1(n_124), .B2(n_386), .ZN(n_385));
   XOR2_X1 i_2 (.A(n_126), .B(n_5742), .Z(n_247));
   XNOR2_X1 i_3 (.A(n_124), .B(n_387), .ZN(n_248));
   INV_X1 i_4 (.A(n_387), .ZN(n_386));
   AOI21_X1 i_5 (.A(n_121), .B1(n_120), .B2(n_454), .ZN(n_387));
   INV_X1 i_6 (.A(n_388), .ZN(n_249));
   AOI21_X1 i_7 (.A(n_123), .B1(n_122), .B2(n_390), .ZN(n_388));
   INV_X1 i_8 (.A(n_389), .ZN(n_250));
   AOI21_X1 i_9 (.A(n_119), .B1(n_118), .B2(n_392), .ZN(n_389));
   XNOR2_X1 i_10 (.A(n_122), .B(n_391), .ZN(n_251));
   INV_X1 i_11 (.A(n_391), .ZN(n_390));
   AOI21_X1 i_12 (.A(n_117), .B1(n_116), .B2(n_393), .ZN(n_391));
   XOR2_X1 i_13 (.A(n_118), .B(n_392), .Z(n_252));
   XOR2_X1 i_14 (.A(n_116), .B(n_393), .Z(n_392));
   XOR2_X1 i_15 (.A(n_460), .B(n_394), .Z(n_393));
   OAI21_X1 i_16 (.A(n_461), .B1(n_484), .B2(n_462), .ZN(n_394));
   INV_X1 i_17 (.A(n_395), .ZN(n_253));
   AOI21_X1 i_18 (.A(n_115), .B1(n_114), .B2(n_397), .ZN(n_395));
   INV_X1 i_19 (.A(n_396), .ZN(n_254));
   AOI21_X1 i_20 (.A(n_109), .B1(n_108), .B2(n_398), .ZN(n_396));
   XOR2_X1 i_21 (.A(n_114), .B(n_397), .Z(n_255));
   XOR2_X1 i_22 (.A(n_112), .B(n_465), .Z(n_397));
   XOR2_X1 i_23 (.A(n_108), .B(n_398), .Z(n_256));
   XNOR2_X1 i_24 (.A(n_106), .B(n_476), .ZN(n_398));
   INV_X1 i_25 (.A(n_399), .ZN(n_257));
   AOI21_X1 i_26 (.A(n_101), .B1(n_100), .B2(n_401), .ZN(n_399));
   INV_X1 i_27 (.A(n_400), .ZN(n_258));
   AOI21_X1 i_28 (.A(n_93), .B1(n_92), .B2(n_403), .ZN(n_400));
   XNOR2_X1 i_29 (.A(n_100), .B(n_402), .ZN(n_259));
   INV_X1 i_30 (.A(n_402), .ZN(n_401));
   AOI21_X1 i_31 (.A(n_91), .B1(n_90), .B2(n_404), .ZN(n_402));
   XOR2_X1 i_32 (.A(n_92), .B(n_403), .Z(n_260));
   XOR2_X1 i_33 (.A(n_90), .B(n_404), .Z(n_403));
   XOR2_X1 i_34 (.A(n_88), .B(n_508), .Z(n_404));
   INV_X1 i_35 (.A(n_405), .ZN(n_261));
   AOI21_X1 i_36 (.A(n_83), .B1(n_82), .B2(n_406), .ZN(n_405));
   XOR2_X1 i_37 (.A(n_82), .B(n_406), .Z(n_262));
   XNOR2_X1 i_38 (.A(n_80), .B(n_535), .ZN(n_406));
   INV_X1 i_39 (.A(n_407), .ZN(n_263));
   AOI21_X1 i_40 (.A(n_71), .B1(n_70), .B2(n_409), .ZN(n_407));
   INV_X1 i_41 (.A(n_408), .ZN(n_264));
   AOI21_X1 i_42 (.A(n_59), .B1(n_58), .B2(n_410), .ZN(n_408));
   XOR2_X1 i_43 (.A(n_70), .B(n_409), .Z(n_265));
   XNOR2_X1 i_44 (.A(n_68), .B(n_561), .ZN(n_409));
   XOR2_X1 i_45 (.A(n_58), .B(n_410), .Z(n_266));
   XNOR2_X1 i_46 (.A(n_56), .B(n_590), .ZN(n_410));
   INV_X1 i_47 (.A(n_411), .ZN(n_267));
   AOI21_X1 i_48 (.A(n_45), .B1(n_44), .B2(n_412), .ZN(n_411));
   XOR2_X1 i_49 (.A(n_44), .B(n_412), .Z(n_268));
   XNOR2_X1 i_50 (.A(n_42), .B(n_624), .ZN(n_412));
   INV_X1 i_51 (.A(n_413), .ZN(n_269));
   AOI21_X1 i_52 (.A(n_29), .B1(n_28), .B2(n_415), .ZN(n_413));
   INV_X1 i_53 (.A(n_414), .ZN(n_270));
   AOI21_X1 i_54 (.A(n_13), .B1(n_12), .B2(n_416), .ZN(n_414));
   XOR2_X1 i_55 (.A(n_28), .B(n_415), .Z(n_271));
   XNOR2_X1 i_56 (.A(n_26), .B(n_671), .ZN(n_415));
   XOR2_X1 i_57 (.A(n_12), .B(n_416), .Z(n_272));
   XNOR2_X1 i_58 (.A(n_10), .B(n_700), .ZN(n_416));
   INV_X1 i_59 (.A(n_417), .ZN(n_5721));
   AOI21_X1 i_60 (.A(n_5718), .B1(n_5717), .B2(n_418), .ZN(n_417));
   XOR2_X1 i_61 (.A(n_5717), .B(n_418), .Z(n_5719));
   XNOR2_X1 i_62 (.A(n_5712), .B(n_748), .ZN(n_418));
   INV_X1 i_63 (.A(n_419), .ZN(n_5635));
   AOI21_X1 i_64 (.A(n_5632), .B1(n_5631), .B2(n_420), .ZN(n_419));
   XOR2_X1 i_65 (.A(n_5631), .B(n_420), .Z(n_5633));
   XNOR2_X1 i_66 (.A(n_5626), .B(n_793), .ZN(n_420));
   INV_X1 i_67 (.A(n_421), .ZN(n_5541));
   AOI21_X1 i_68 (.A(n_5538), .B1(n_5537), .B2(n_422), .ZN(n_421));
   XOR2_X1 i_69 (.A(n_5537), .B(n_422), .Z(n_5539));
   XNOR2_X1 i_70 (.A(n_5532), .B(n_840), .ZN(n_422));
   INV_X1 i_71 (.A(n_423), .ZN(n_5442));
   AOI21_X1 i_72 (.A(n_5439), .B1(n_5438), .B2(n_424), .ZN(n_423));
   XOR2_X1 i_73 (.A(n_5438), .B(n_424), .Z(n_5440));
   XNOR2_X1 i_74 (.A(n_5433), .B(n_897), .ZN(n_424));
   INV_X1 i_75 (.A(n_425), .ZN(n_5339));
   AOI21_X1 i_76 (.A(n_5336), .B1(n_5335), .B2(n_426), .ZN(n_425));
   XOR2_X1 i_77 (.A(n_5335), .B(n_426), .Z(n_5337));
   XNOR2_X1 i_78 (.A(n_5330), .B(n_954), .ZN(n_426));
   INV_X1 i_79 (.A(n_427), .ZN(n_5228));
   AOI21_X1 i_80 (.A(n_5225), .B1(n_5224), .B2(n_428), .ZN(n_427));
   XOR2_X1 i_81 (.A(n_5224), .B(n_428), .Z(n_5226));
   XNOR2_X1 i_82 (.A(n_5219), .B(n_1014), .ZN(n_428));
   INV_X1 i_83 (.A(n_429), .ZN(n_5112));
   AOI21_X1 i_84 (.A(n_5109), .B1(n_5108), .B2(n_430), .ZN(n_429));
   XOR2_X1 i_85 (.A(n_5108), .B(n_430), .Z(n_5110));
   XOR2_X1 i_86 (.A(n_5103), .B(n_1109), .Z(n_430));
   INV_X1 i_87 (.A(n_431), .ZN(n_4992));
   AOI21_X1 i_88 (.A(n_4989), .B1(n_4988), .B2(n_432), .ZN(n_431));
   XOR2_X1 i_89 (.A(n_4988), .B(n_432), .Z(n_4990));
   XNOR2_X1 i_90 (.A(n_4983), .B(n_1218), .ZN(n_432));
   INV_X1 i_91 (.A(n_433), .ZN(n_4864));
   AOI21_X1 i_92 (.A(n_4861), .B1(n_4860), .B2(n_434), .ZN(n_433));
   XOR2_X1 i_93 (.A(n_4860), .B(n_434), .Z(n_4862));
   XNOR2_X1 i_94 (.A(n_4855), .B(n_1336), .ZN(n_434));
   INV_X1 i_95 (.A(n_435), .ZN(n_4731));
   AOI21_X1 i_96 (.A(n_4728), .B1(n_4727), .B2(n_436), .ZN(n_435));
   XOR2_X1 i_97 (.A(n_4727), .B(n_436), .Z(n_4729));
   XNOR2_X1 i_98 (.A(n_4722), .B(n_1464), .ZN(n_436));
   INV_X1 i_99 (.A(n_437), .ZN(n_4594));
   AOI21_X1 i_100 (.A(n_4591), .B1(n_4590), .B2(n_438), .ZN(n_437));
   XOR2_X1 i_101 (.A(n_4590), .B(n_438), .Z(n_4592));
   XNOR2_X1 i_102 (.A(n_4585), .B(n_1592), .ZN(n_438));
   INV_X1 i_103 (.A(n_439), .ZN(n_4449));
   AOI21_X1 i_104 (.A(n_4446), .B1(n_4445), .B2(n_440), .ZN(n_439));
   XOR2_X1 i_105 (.A(n_4445), .B(n_440), .Z(n_4447));
   XNOR2_X1 i_106 (.A(n_4440), .B(n_1725), .ZN(n_440));
   INV_X1 i_107 (.A(n_441), .ZN(n_4299));
   AOI21_X1 i_108 (.A(n_4296), .B1(n_4295), .B2(n_443), .ZN(n_441));
   INV_X1 i_109 (.A(n_442), .ZN(n_4145));
   AOI21_X1 i_110 (.A(n_4142), .B1(n_4141), .B2(n_444), .ZN(n_442));
   XOR2_X1 i_111 (.A(n_4295), .B(n_443), .Z(n_4297));
   XOR2_X1 i_112 (.A(n_4290), .B(n_1868), .Z(n_443));
   XOR2_X1 i_113 (.A(n_4141), .B(n_444), .Z(n_4143));
   XNOR2_X1 i_114 (.A(n_4136), .B(n_2018), .ZN(n_444));
   INV_X1 i_115 (.A(n_445), .ZN(n_3983));
   AOI21_X1 i_116 (.A(n_3980), .B1(n_3979), .B2(n_446), .ZN(n_445));
   XOR2_X1 i_117 (.A(n_3979), .B(n_446), .Z(n_3981));
   XNOR2_X1 i_118 (.A(n_3974), .B(n_2155), .ZN(n_446));
   INV_X1 i_119 (.A(n_448), .ZN(n_3816));
   AOI21_X1 i_120 (.A(n_3813), .B1(n_3812), .B2(n_449), .ZN(n_448));
   XNOR2_X1 i_121 (.A(n_3812), .B(n_450), .ZN(n_3814));
   INV_X1 i_122 (.A(n_450), .ZN(n_449));
   AOI21_X1 i_123 (.A(n_3641), .B1(n_3640), .B2(n_2644), .ZN(n_450));
   XOR2_X1 i_124 (.A(n_2706), .B(n_3509), .Z(n_2708));
   XOR2_X1 i_125 (.A(n_2083), .B(n_4205), .Z(n_2085));
   XOR2_X1 i_126 (.A(n_1778), .B(n_4563), .Z(n_1780));
   XOR2_X1 i_127 (.A(n_1689), .B(n_4655), .Z(n_1691));
   XOR2_X1 i_128 (.A(n_1604), .B(n_4762), .Z(n_1606));
   XOR2_X1 i_129 (.A(n_1524), .B(n_4873), .Z(n_1526));
   XNOR2_X1 i_130 (.A(n_1452), .B(n_4951), .ZN(n_1454));
   XOR2_X1 i_131 (.A(n_1384), .B(n_4956), .Z(n_1386));
   XOR2_X1 i_132 (.A(n_1321), .B(n_5118), .Z(n_1323));
   XOR2_X1 i_133 (.A(n_1266), .B(n_5159), .Z(n_1268));
   XOR2_X1 i_134 (.A(n_1215), .B(n_5238), .Z(n_1217));
   XOR2_X1 i_135 (.A(n_1137), .B(n_1169), .Z(n_1171));
   XOR2_X1 i_136 (.A(n_1103), .B(n_1131), .Z(n_1133));
   XOR2_X1 i_137 (.A(n_1097), .B(n_5368), .Z(n_1099));
   XOR2_X1 i_138 (.A(n_1068), .B(n_5426), .Z(n_1070));
   XOR2_X1 i_139 (.A(n_5465), .B(n_451), .Z(n_1039));
   NAND2_X1 i_140 (.A1(n_5470), .A2(n_5466), .ZN(n_451));
   XOR2_X1 i_141 (.A(n_5480), .B(n_452), .Z(n_1029));
   NAND2_X1 i_142 (.A1(n_5483), .A2(n_5481), .ZN(n_452));
   OAI22_X1 i_143 (.A1(n_5495), .A2(n_5477), .B1(n_5496), .B2(n_5478), .ZN(
      n_1034));
   NAND2_X1 i_144 (.A1(inputB[30]), .A2(inputA[31]), .ZN(n_991));
   NAND2_X1 i_145 (.A1(inputB[31]), .A2(inputA[30]), .ZN(n_1022));
   XOR2_X1 i_146 (.A(n_5745), .B(n_5743), .Z(n_273));
   INV_X1 i_147 (.A(n_453), .ZN(n_274));
   AOI22_X1 i_148 (.A1(n_5748), .A2(n_462), .B1(n_458), .B2(n_457), .ZN(n_453));
   XNOR2_X1 i_149 (.A(n_120), .B(n_455), .ZN(n_275));
   INV_X1 i_150 (.A(n_455), .ZN(n_454));
   AOI21_X1 i_151 (.A(n_456), .B1(n_473), .B2(n_470), .ZN(n_455));
   AOI21_X1 i_152 (.A(n_471), .B1(n_472), .B2(n_469), .ZN(n_456));
   XOR2_X1 i_153 (.A(n_458), .B(n_457), .Z(n_276));
   NAND2_X1 i_154 (.A1(inputB[31]), .A2(inputA[28]), .ZN(n_457));
   AOI21_X1 i_155 (.A(n_459), .B1(n_5748), .B2(n_462), .ZN(n_458));
   AOI22_X1 i_156 (.A1(inputB[30]), .A2(inputA[29]), .B1(inputB[29]), .B2(
      inputA[30]), .ZN(n_459));
   AOI22_X1 i_157 (.A1(n_485), .A2(n_463), .B1(n_461), .B2(n_460), .ZN(n_277));
   AND2_X1 i_158 (.A1(inputB[31]), .A2(inputA[27]), .ZN(n_460));
   NAND2_X1 i_159 (.A1(n_484), .A2(n_462), .ZN(n_461));
   INV_X1 i_160 (.A(n_463), .ZN(n_462));
   NAND2_X1 i_161 (.A1(inputB[29]), .A2(inputA[29]), .ZN(n_463));
   NAND2_X1 i_162 (.A1(inputB[28]), .A2(inputA[31]), .ZN(n_927));
   INV_X1 i_163 (.A(n_464), .ZN(n_278));
   AOI21_X1 i_164 (.A(n_113), .B1(n_112), .B2(n_465), .ZN(n_464));
   XNOR2_X1 i_165 (.A(n_110), .B(n_468), .ZN(n_465));
   INV_X1 i_166 (.A(n_466), .ZN(n_279));
   AOI21_X1 i_167 (.A(n_111), .B1(n_110), .B2(n_467), .ZN(n_466));
   INV_X1 i_168 (.A(n_468), .ZN(n_467));
   AOI21_X1 i_169 (.A(n_103), .B1(n_102), .B2(n_499), .ZN(n_468));
   XOR2_X1 i_170 (.A(n_473), .B(n_469), .Z(n_280));
   XNOR2_X1 i_171 (.A(n_471), .B(n_470), .ZN(n_469));
   NAND2_X1 i_172 (.A1(inputB[27]), .A2(inputA[31]), .ZN(n_470));
   NAND2_X1 i_173 (.A1(inputB[28]), .A2(inputA[30]), .ZN(n_471));
   INV_X1 i_174 (.A(n_473), .ZN(n_472));
   AOI21_X1 i_175 (.A(n_488), .B1(n_489), .B2(n_486), .ZN(n_473));
   AOI21_X1 i_176 (.A(n_482), .B1(n_483), .B2(n_478), .ZN(n_281));
   INV_X1 i_177 (.A(n_474), .ZN(n_282));
   AOI21_X1 i_178 (.A(n_107), .B1(n_106), .B2(n_475), .ZN(n_474));
   INV_X1 i_179 (.A(n_476), .ZN(n_475));
   AOI21_X1 i_180 (.A(n_97), .B1(n_96), .B2(n_509), .ZN(n_476));
   INV_X1 i_181 (.A(n_477), .ZN(n_283));
   AOI21_X1 i_182 (.A(n_105), .B1(n_104), .B2(n_492), .ZN(n_477));
   XNOR2_X1 i_183 (.A(n_480), .B(n_479), .ZN(n_284));
   INV_X1 i_184 (.A(n_479), .ZN(n_478));
   NAND2_X1 i_185 (.A1(inputB[31]), .A2(inputA[26]), .ZN(n_479));
   NAND2_X1 i_186 (.A1(n_483), .A2(n_481), .ZN(n_480));
   INV_X1 i_187 (.A(n_482), .ZN(n_481));
   AOI22_X1 i_188 (.A1(inputB[30]), .A2(inputA[27]), .B1(inputB[29]), .B2(
      inputA[28]), .ZN(n_482));
   NAND2_X1 i_189 (.A1(n_498), .A2(n_484), .ZN(n_483));
   INV_X1 i_190 (.A(n_485), .ZN(n_484));
   NAND2_X1 i_191 (.A1(inputB[30]), .A2(inputA[28]), .ZN(n_485));
   XNOR2_X1 i_192 (.A(n_487), .B(n_486), .ZN(n_285));
   NAND2_X1 i_193 (.A1(inputB[28]), .A2(inputA[29]), .ZN(n_486));
   NOR2_X1 i_194 (.A1(n_490), .A2(n_488), .ZN(n_487));
   AND3_X1 i_195 (.A1(inputB[26]), .A2(inputA[31]), .A3(n_503), .ZN(n_488));
   INV_X1 i_196 (.A(n_490), .ZN(n_489));
   AOI21_X1 i_197 (.A(n_503), .B1(inputB[26]), .B2(inputA[31]), .ZN(n_490));
   AOI21_X1 i_198 (.A(n_497), .B1(n_496), .B2(n_493), .ZN(n_286));
   OAI22_X1 i_199 (.A1(n_525), .A2(n_503), .B1(n_505), .B2(n_501), .ZN(n_287));
   INV_X1 i_200 (.A(n_491), .ZN(n_288));
   AOI21_X1 i_201 (.A(n_99), .B1(n_98), .B2(n_506), .ZN(n_491));
   XOR2_X1 i_202 (.A(n_104), .B(n_492), .Z(n_289));
   XNOR2_X1 i_203 (.A(n_494), .B(n_493), .ZN(n_492));
   AND2_X1 i_204 (.A1(inputB[31]), .A2(inputA[25]), .ZN(n_493));
   NOR2_X1 i_205 (.A1(n_497), .A2(n_495), .ZN(n_494));
   INV_X1 i_206 (.A(n_496), .ZN(n_495));
   NAND3_X1 i_207 (.A1(inputB[30]), .A2(inputA[26]), .A3(n_498), .ZN(n_496));
   AOI21_X1 i_208 (.A(n_498), .B1(inputB[30]), .B2(inputA[26]), .ZN(n_497));
   AND2_X1 i_209 (.A1(inputB[29]), .A2(inputA[27]), .ZN(n_498));
   XOR2_X1 i_210 (.A(n_102), .B(n_499), .Z(n_290));
   OAI21_X1 i_211 (.A(n_514), .B1(n_515), .B2(n_510), .ZN(n_499));
   INV_X1 i_212 (.A(n_500), .ZN(n_291));
   AOI21_X1 i_213 (.A(n_95), .B1(n_94), .B2(n_517), .ZN(n_500));
   XOR2_X1 i_214 (.A(n_502), .B(n_501), .Z(n_292));
   NAND2_X1 i_215 (.A1(inputB[28]), .A2(inputA[28]), .ZN(n_501));
   OAI21_X1 i_216 (.A(n_504), .B1(n_525), .B2(n_503), .ZN(n_502));
   NAND2_X1 i_217 (.A1(inputB[27]), .A2(inputA[30]), .ZN(n_503));
   INV_X1 i_218 (.A(n_505), .ZN(n_504));
   AOI22_X1 i_219 (.A1(inputB[27]), .A2(inputA[29]), .B1(inputB[26]), .B2(
      inputA[30]), .ZN(n_505));
   AOI21_X1 i_220 (.A(n_531), .B1(n_530), .B2(n_526), .ZN(n_293));
   AOI22_X1 i_221 (.A1(n_545), .A2(n_525), .B1(n_523), .B2(n_521), .ZN(n_294));
   NAND2_X1 i_222 (.A1(inputB[25]), .A2(inputA[31]), .ZN(n_831));
   XNOR2_X1 i_223 (.A(n_98), .B(n_507), .ZN(n_295));
   INV_X1 i_224 (.A(n_507), .ZN(n_506));
   AOI21_X1 i_225 (.A(n_89), .B1(n_88), .B2(n_508), .ZN(n_507));
   XOR2_X1 i_226 (.A(n_84), .B(n_519), .Z(n_508));
   XOR2_X1 i_227 (.A(n_96), .B(n_509), .Z(n_296));
   XOR2_X1 i_228 (.A(n_512), .B(n_511), .Z(n_509));
   INV_X1 i_229 (.A(n_511), .ZN(n_510));
   NAND2_X1 i_230 (.A1(inputB[31]), .A2(inputA[24]), .ZN(n_511));
   NOR2_X1 i_231 (.A1(n_515), .A2(n_513), .ZN(n_512));
   INV_X1 i_232 (.A(n_514), .ZN(n_513));
   NAND3_X1 i_233 (.A1(inputB[29]), .A2(inputA[26]), .A3(n_551), .ZN(n_514));
   AOI21_X1 i_234 (.A(n_551), .B1(inputB[29]), .B2(inputA[26]), .ZN(n_515));
   INV_X1 i_235 (.A(n_516), .ZN(n_297));
   AOI21_X1 i_236 (.A(n_87), .B1(n_86), .B2(n_537), .ZN(n_516));
   XNOR2_X1 i_237 (.A(n_94), .B(n_518), .ZN(n_298));
   INV_X1 i_238 (.A(n_518), .ZN(n_517));
   AOI21_X1 i_239 (.A(n_85), .B1(n_84), .B2(n_519), .ZN(n_518));
   NAND2_X1 i_240 (.A1(n_570), .A2(n_520), .ZN(n_519));
   NAND2_X1 i_241 (.A1(n_569), .A2(n_567), .ZN(n_520));
   XOR2_X1 i_242 (.A(n_522), .B(n_521), .Z(n_299));
   NAND2_X1 i_243 (.A1(inputB[28]), .A2(inputA[27]), .ZN(n_521));
   OAI21_X1 i_244 (.A(n_523), .B1(n_544), .B2(n_524), .ZN(n_522));
   NAND2_X1 i_245 (.A1(n_544), .A2(n_524), .ZN(n_523));
   INV_X1 i_246 (.A(n_525), .ZN(n_524));
   NAND2_X1 i_247 (.A1(inputB[26]), .A2(inputA[29]), .ZN(n_525));
   XOR2_X1 i_248 (.A(n_528), .B(n_527), .Z(n_300));
   INV_X1 i_249 (.A(n_527), .ZN(n_526));
   AOI21_X1 i_250 (.A(n_554), .B1(n_556), .B2(n_552), .ZN(n_527));
   NOR2_X1 i_251 (.A1(n_531), .A2(n_529), .ZN(n_528));
   INV_X1 i_252 (.A(n_530), .ZN(n_529));
   OAI211_X1 i_253 (.A(inputB[25]), .B(inputA[30]), .C1(n_5767), .C2(n_5753), 
      .ZN(n_530));
   AOI211_X1 i_254 (.A(n_5767), .B(n_5753), .C1(inputB[25]), .C2(inputA[30]), 
      .ZN(n_531));
   INV_X1 i_255 (.A(n_532), .ZN(n_301));
   AOI22_X1 i_256 (.A1(n_571), .A2(n_551), .B1(n_549), .B2(n_548), .ZN(n_532));
   OAI21_X1 i_257 (.A(n_542), .B1(n_541), .B2(n_538), .ZN(n_302));
   INV_X1 i_258 (.A(n_533), .ZN(n_303));
   AOI21_X1 i_259 (.A(n_81), .B1(n_80), .B2(n_534), .ZN(n_533));
   INV_X1 i_260 (.A(n_535), .ZN(n_534));
   AOI21_X1 i_261 (.A(n_67), .B1(n_66), .B2(n_591), .ZN(n_535));
   INV_X1 i_262 (.A(n_536), .ZN(n_304));
   AOI21_X1 i_263 (.A(n_79), .B1(n_78), .B2(n_562), .ZN(n_536));
   XOR2_X1 i_264 (.A(n_86), .B(n_537), .Z(n_305));
   XOR2_X1 i_265 (.A(n_539), .B(n_538), .Z(n_537));
   NAND2_X1 i_266 (.A1(inputB[28]), .A2(inputA[26]), .ZN(n_538));
   NAND2_X1 i_267 (.A1(n_542), .A2(n_540), .ZN(n_539));
   INV_X1 i_268 (.A(n_541), .ZN(n_540));
   AOI22_X1 i_269 (.A1(inputB[27]), .A2(inputA[27]), .B1(inputB[26]), .B2(
      inputA[28]), .ZN(n_541));
   NAND2_X1 i_270 (.A1(n_579), .A2(n_544), .ZN(n_542));
   INV_X1 i_271 (.A(n_545), .ZN(n_544));
   NAND2_X1 i_272 (.A1(inputB[27]), .A2(inputA[28]), .ZN(n_545));
   INV_X1 i_273 (.A(n_546), .ZN(n_306));
   AOI21_X1 i_274 (.A(n_77), .B1(n_76), .B2(n_566), .ZN(n_546));
   INV_X1 i_275 (.A(n_547), .ZN(n_307));
   AOI21_X1 i_276 (.A(n_75), .B1(n_74), .B2(n_563), .ZN(n_547));
   XOR2_X1 i_277 (.A(n_549), .B(n_548), .Z(n_308));
   NAND2_X1 i_278 (.A1(inputB[31]), .A2(inputA[23]), .ZN(n_548));
   AOI21_X1 i_279 (.A(n_550), .B1(n_571), .B2(n_551), .ZN(n_549));
   AOI22_X1 i_280 (.A1(inputB[30]), .A2(inputA[24]), .B1(inputB[29]), .B2(
      inputA[25]), .ZN(n_550));
   AND2_X1 i_281 (.A1(inputB[30]), .A2(inputA[25]), .ZN(n_551));
   XNOR2_X1 i_282 (.A(n_553), .B(n_552), .ZN(n_309));
   NAND2_X1 i_283 (.A1(inputB[25]), .A2(inputA[29]), .ZN(n_552));
   NOR2_X1 i_284 (.A1(n_555), .A2(n_554), .ZN(n_553));
   AOI21_X1 i_285 (.A(n_557), .B1(inputB[24]), .B2(inputA[30]), .ZN(n_554));
   INV_X1 i_286 (.A(n_556), .ZN(n_555));
   NAND3_X1 i_287 (.A1(inputB[24]), .A2(inputA[30]), .A3(n_557), .ZN(n_556));
   NAND2_X1 i_288 (.A1(inputB[23]), .A2(inputA[31]), .ZN(n_557));
   INV_X1 i_289 (.A(n_558), .ZN(n_310));
   AOI21_X1 i_290 (.A(n_73), .B1(n_72), .B2(n_575), .ZN(n_558));
   AOI22_X1 i_291 (.A1(n_613), .A2(n_580), .B1(n_578), .B2(n_576), .ZN(n_311));
   OAI21_X1 i_292 (.A(n_583), .B1(n_585), .B2(n_581), .ZN(n_312));
   INV_X1 i_293 (.A(n_559), .ZN(n_313));
   AOI21_X1 i_294 (.A(n_69), .B1(n_68), .B2(n_560), .ZN(n_559));
   INV_X1 i_295 (.A(n_561), .ZN(n_560));
   AOI21_X1 i_296 (.A(n_55), .B1(n_54), .B2(n_625), .ZN(n_561));
   XOR2_X1 i_297 (.A(n_78), .B(n_562), .Z(n_314));
   XNOR2_X1 i_298 (.A(n_74), .B(n_564), .ZN(n_562));
   INV_X1 i_299 (.A(n_564), .ZN(n_563));
   AOI21_X1 i_300 (.A(n_565), .B1(n_618), .B2(n_617), .ZN(n_564));
   AOI21_X1 i_301 (.A(n_645), .B1(n_619), .B2(n_616), .ZN(n_565));
   XOR2_X1 i_302 (.A(n_76), .B(n_566), .Z(n_315));
   XOR2_X1 i_303 (.A(n_568), .B(n_567), .Z(n_566));
   NAND2_X1 i_304 (.A1(inputB[31]), .A2(inputA[22]), .ZN(n_567));
   AND2_X1 i_305 (.A1(n_570), .A2(n_569), .ZN(n_568));
   NAND2_X1 i_306 (.A1(n_608), .A2(n_572), .ZN(n_569));
   NAND2_X1 i_307 (.A1(n_607), .A2(n_571), .ZN(n_570));
   INV_X1 i_308 (.A(n_572), .ZN(n_571));
   NAND2_X1 i_309 (.A1(inputB[29]), .A2(inputA[24]), .ZN(n_572));
   INV_X1 i_310 (.A(n_573), .ZN(n_316));
   AOI21_X1 i_311 (.A(n_65), .B1(n_64), .B2(n_600), .ZN(n_573));
   INV_X1 i_312 (.A(n_574), .ZN(n_317));
   AOI21_X1 i_313 (.A(n_63), .B1(n_62), .B2(n_593), .ZN(n_574));
   XOR2_X1 i_314 (.A(n_72), .B(n_575), .Z(n_318));
   OAI21_X1 i_315 (.A(n_611), .B1(n_615), .B2(n_609), .ZN(n_575));
   XOR2_X1 i_316 (.A(n_577), .B(n_576), .Z(n_319));
   NAND2_X1 i_317 (.A1(inputB[28]), .A2(inputA[25]), .ZN(n_576));
   OAI21_X1 i_318 (.A(n_578), .B1(n_612), .B2(n_579), .ZN(n_577));
   NAND2_X1 i_319 (.A1(n_612), .A2(n_579), .ZN(n_578));
   INV_X1 i_320 (.A(n_580), .ZN(n_579));
   NAND2_X1 i_321 (.A1(inputB[26]), .A2(inputA[27]), .ZN(n_580));
   XOR2_X1 i_322 (.A(n_582), .B(n_581), .Z(n_320));
   NAND2_X1 i_323 (.A1(inputB[25]), .A2(inputA[28]), .ZN(n_581));
   NAND2_X1 i_324 (.A1(n_584), .A2(n_583), .ZN(n_582));
   NAND3_X1 i_325 (.A1(inputB[23]), .A2(inputA[30]), .A3(n_599), .ZN(n_583));
   INV_X1 i_326 (.A(n_585), .ZN(n_584));
   AOI21_X1 i_327 (.A(n_599), .B1(inputB[23]), .B2(inputA[30]), .ZN(n_585));
   INV_X1 i_328 (.A(n_586), .ZN(n_321));
   AOI21_X1 i_329 (.A(n_61), .B1(n_60), .B2(n_601), .ZN(n_586));
   NOR2_X1 i_330 (.A1(n_606), .A2(n_587), .ZN(n_322));
   AOI21_X1 i_331 (.A(n_604), .B1(n_635), .B2(n_607), .ZN(n_587));
   OAI21_X1 i_332 (.A(n_598), .B1(n_597), .B2(n_594), .ZN(n_323));
   NAND2_X1 i_333 (.A1(inputB[22]), .A2(inputA[31]), .ZN(n_735));
   INV_X1 i_334 (.A(n_588), .ZN(n_324));
   AOI21_X1 i_335 (.A(n_57), .B1(n_56), .B2(n_589), .ZN(n_588));
   INV_X1 i_336 (.A(n_590), .ZN(n_589));
   AOI21_X1 i_337 (.A(n_41), .B1(n_40), .B2(n_660), .ZN(n_590));
   XNOR2_X1 i_338 (.A(n_66), .B(n_592), .ZN(n_325));
   INV_X1 i_339 (.A(n_592), .ZN(n_591));
   AOI21_X1 i_340 (.A(n_53), .B1(n_52), .B2(n_627), .ZN(n_592));
   XOR2_X1 i_341 (.A(n_62), .B(n_593), .Z(n_326));
   XOR2_X1 i_342 (.A(n_595), .B(n_594), .Z(n_593));
   NAND2_X1 i_343 (.A1(inputB[25]), .A2(inputA[27]), .ZN(n_594));
   NAND2_X1 i_344 (.A1(n_598), .A2(n_596), .ZN(n_595));
   INV_X1 i_345 (.A(n_597), .ZN(n_596));
   AOI22_X1 i_346 (.A1(inputB[24]), .A2(inputA[28]), .B1(inputB[23]), .B2(
      inputA[29]), .ZN(n_597));
   NAND2_X1 i_347 (.A1(n_657), .A2(n_599), .ZN(n_598));
   NOR2_X1 i_348 (.A1(n_5767), .A2(n_5750), .ZN(n_599));
   XOR2_X1 i_349 (.A(n_64), .B(n_600), .Z(n_327));
   XOR2_X1 i_350 (.A(n_60), .B(n_601), .Z(n_600));
   NAND2_X1 i_351 (.A1(n_634), .A2(n_630), .ZN(n_601));
   INV_X1 i_352 (.A(n_602), .ZN(n_328));
   AOI21_X1 i_353 (.A(n_49), .B1(n_48), .B2(n_638), .ZN(n_602));
   INV_X1 i_354 (.A(n_603), .ZN(n_329));
   AOI21_X1 i_355 (.A(n_51), .B1(n_50), .B2(n_629), .ZN(n_603));
   XOR2_X1 i_356 (.A(n_605), .B(n_604), .Z(n_330));
   NAND2_X1 i_357 (.A1(inputB[31]), .A2(inputA[21]), .ZN(n_604));
   AOI21_X1 i_358 (.A(n_606), .B1(n_635), .B2(n_607), .ZN(n_605));
   AOI22_X1 i_359 (.A1(inputB[30]), .A2(inputA[22]), .B1(inputB[29]), .B2(
      inputA[23]), .ZN(n_606));
   INV_X1 i_360 (.A(n_608), .ZN(n_607));
   NAND2_X1 i_361 (.A1(inputB[30]), .A2(inputA[23]), .ZN(n_608));
   XOR2_X1 i_362 (.A(n_610), .B(n_609), .Z(n_331));
   NAND2_X1 i_363 (.A1(inputB[28]), .A2(inputA[24]), .ZN(n_609));
   NAND2_X1 i_364 (.A1(n_614), .A2(n_611), .ZN(n_610));
   NAND3_X1 i_365 (.A1(inputB[26]), .A2(inputA[25]), .A3(n_612), .ZN(n_611));
   INV_X1 i_366 (.A(n_613), .ZN(n_612));
   NAND2_X1 i_367 (.A1(inputB[27]), .A2(inputA[26]), .ZN(n_613));
   INV_X1 i_368 (.A(n_615), .ZN(n_614));
   AOI22_X1 i_369 (.A1(inputB[27]), .A2(inputA[25]), .B1(inputB[26]), .B2(
      inputA[26]), .ZN(n_615));
   XOR2_X1 i_370 (.A(n_618), .B(n_616), .Z(n_332));
   XNOR2_X1 i_371 (.A(n_645), .B(n_617), .ZN(n_616));
   NAND2_X1 i_372 (.A1(inputB[21]), .A2(inputA[31]), .ZN(n_617));
   INV_X1 i_373 (.A(n_619), .ZN(n_618));
   AOI21_X1 i_374 (.A(n_644), .B1(n_642), .B2(n_640), .ZN(n_619));
   INV_X1 i_375 (.A(n_620), .ZN(n_333));
   AOI21_X1 i_376 (.A(n_47), .B1(n_46), .B2(n_646), .ZN(n_620));
   OAI21_X1 i_377 (.A(n_650), .B1(n_652), .B2(n_648), .ZN(n_334));
   NAND2_X1 i_378 (.A1(n_656), .A2(n_621), .ZN(n_335));
   NAND2_X1 i_379 (.A1(n_655), .A2(n_653), .ZN(n_621));
   INV_X1 i_380 (.A(n_622), .ZN(n_336));
   AOI21_X1 i_381 (.A(n_43), .B1(n_42), .B2(n_623), .ZN(n_622));
   INV_X1 i_382 (.A(n_624), .ZN(n_623));
   AOI21_X1 i_383 (.A(n_25), .B1(n_24), .B2(n_701), .ZN(n_624));
   XNOR2_X1 i_384 (.A(n_54), .B(n_626), .ZN(n_337));
   INV_X1 i_385 (.A(n_626), .ZN(n_625));
   AOI21_X1 i_386 (.A(n_37), .B1(n_36), .B2(n_675), .ZN(n_626));
   XNOR2_X1 i_387 (.A(n_52), .B(n_628), .ZN(n_338));
   INV_X1 i_388 (.A(n_628), .ZN(n_627));
   AOI21_X1 i_389 (.A(n_35), .B1(n_34), .B2(n_661), .ZN(n_628));
   XOR2_X1 i_390 (.A(n_50), .B(n_629), .Z(n_339));
   XNOR2_X1 i_391 (.A(n_632), .B(n_631), .ZN(n_629));
   NAND2_X1 i_392 (.A1(n_633), .A2(n_631), .ZN(n_630));
   NAND2_X1 i_393 (.A1(inputB[31]), .A2(inputA[20]), .ZN(n_631));
   NAND2_X1 i_394 (.A1(n_634), .A2(n_633), .ZN(n_632));
   NAND2_X1 i_395 (.A1(n_685), .A2(n_636), .ZN(n_633));
   NAND2_X1 i_396 (.A1(n_684), .A2(n_635), .ZN(n_634));
   INV_X1 i_397 (.A(n_636), .ZN(n_635));
   NAND2_X1 i_398 (.A1(inputB[29]), .A2(inputA[22]), .ZN(n_636));
   INV_X1 i_399 (.A(n_637), .ZN(n_340));
   AOI21_X1 i_400 (.A(n_39), .B1(n_38), .B2(n_672), .ZN(n_637));
   XOR2_X1 i_401 (.A(n_48), .B(n_638), .Z(n_341));
   XOR2_X1 i_402 (.A(n_641), .B(n_640), .Z(n_638));
   NAND2_X1 i_403 (.A1(inputB[20]), .A2(inputA[31]), .ZN(n_640));
   NOR2_X1 i_404 (.A1(n_644), .A2(n_643), .ZN(n_641));
   INV_X1 i_405 (.A(n_643), .ZN(n_642));
   AOI22_X1 i_406 (.A1(inputB[21]), .A2(inputA[30]), .B1(inputB[22]), .B2(
      inputA[29]), .ZN(n_643));
   NOR2_X1 i_407 (.A1(n_742), .A2(n_645), .ZN(n_644));
   NAND2_X1 i_408 (.A1(inputB[22]), .A2(inputA[30]), .ZN(n_645));
   XOR2_X1 i_409 (.A(n_46), .B(n_646), .Z(n_342));
   AOI22_X1 i_410 (.A1(n_721), .A2(n_692), .B1(n_690), .B2(n_688), .ZN(n_646));
   INV_X1 i_411 (.A(n_647), .ZN(n_343));
   AOI21_X1 i_412 (.A(n_33), .B1(n_32), .B2(n_676), .ZN(n_647));
   XOR2_X1 i_413 (.A(n_649), .B(n_648), .Z(n_344));
   NAND2_X1 i_414 (.A1(inputB[28]), .A2(inputA[23]), .ZN(n_648));
   NAND2_X1 i_415 (.A1(n_651), .A2(n_650), .ZN(n_649));
   NAND3_X1 i_416 (.A1(inputB[27]), .A2(inputA[25]), .A3(n_691), .ZN(n_650));
   INV_X1 i_417 (.A(n_652), .ZN(n_651));
   AOI22_X1 i_418 (.A1(inputB[27]), .A2(inputA[24]), .B1(inputB[26]), .B2(
      inputA[25]), .ZN(n_652));
   XOR2_X1 i_419 (.A(n_654), .B(n_653), .Z(n_345));
   AND2_X1 i_420 (.A1(inputB[25]), .A2(inputA[26]), .ZN(n_653));
   AND2_X1 i_421 (.A1(n_656), .A2(n_655), .ZN(n_654));
   NAND2_X1 i_422 (.A1(n_668), .A2(n_658), .ZN(n_655));
   NAND2_X1 i_423 (.A1(n_667), .A2(n_657), .ZN(n_656));
   INV_X1 i_424 (.A(n_658), .ZN(n_657));
   NAND2_X1 i_425 (.A1(inputB[23]), .A2(inputA[28]), .ZN(n_658));
   INV_X1 i_426 (.A(n_659), .ZN(n_346));
   AOI21_X1 i_427 (.A(n_31), .B1(n_30), .B2(n_680), .ZN(n_659));
   AOI21_X1 i_428 (.A(n_686), .B1(n_687), .B2(n_683), .ZN(n_347));
   OAI21_X1 i_429 (.A(n_666), .B1(n_665), .B2(n_662), .ZN(n_348));
   OAI21_X1 i_430 (.A(n_697), .B1(n_695), .B2(n_693), .ZN(n_349));
   XOR2_X1 i_431 (.A(n_40), .B(n_660), .Z(n_350));
   XOR2_X1 i_432 (.A(n_34), .B(n_661), .Z(n_660));
   XOR2_X1 i_433 (.A(n_663), .B(n_662), .Z(n_661));
   NAND2_X1 i_434 (.A1(inputB[25]), .A2(inputA[25]), .ZN(n_662));
   NAND2_X1 i_435 (.A1(n_666), .A2(n_664), .ZN(n_663));
   INV_X1 i_436 (.A(n_665), .ZN(n_664));
   AOI22_X1 i_437 (.A1(inputB[24]), .A2(inputA[26]), .B1(inputB[23]), .B2(
      inputA[27]), .ZN(n_665));
   NAND2_X1 i_438 (.A1(n_737), .A2(n_667), .ZN(n_666));
   INV_X1 i_439 (.A(n_668), .ZN(n_667));
   NAND2_X1 i_440 (.A1(inputB[24]), .A2(inputA[27]), .ZN(n_668));
   INV_X1 i_441 (.A(n_669), .ZN(n_351));
   AOI21_X1 i_442 (.A(n_27), .B1(n_26), .B2(n_670), .ZN(n_669));
   INV_X1 i_443 (.A(n_671), .ZN(n_670));
   AOI21_X1 i_444 (.A(n_9), .B1(n_8), .B2(n_749), .ZN(n_671));
   XNOR2_X1 i_445 (.A(n_38), .B(n_673), .ZN(n_352));
   INV_X1 i_446 (.A(n_673), .ZN(n_672));
   AOI21_X1 i_447 (.A(n_17), .B1(n_16), .B2(n_706), .ZN(n_673));
   INV_X1 i_448 (.A(n_674), .ZN(n_353));
   AOI21_X1 i_449 (.A(n_23), .B1(n_22), .B2(n_705), .ZN(n_674));
   XOR2_X1 i_450 (.A(n_36), .B(n_675), .Z(n_354));
   XNOR2_X1 i_451 (.A(n_32), .B(n_677), .ZN(n_675));
   INV_X1 i_452 (.A(n_677), .ZN(n_676));
   AOI21_X1 i_453 (.A(n_15), .B1(n_14), .B2(n_703), .ZN(n_677));
   INV_X1 i_454 (.A(n_678), .ZN(n_355));
   AOI21_X1 i_455 (.A(n_21), .B1(n_20), .B2(n_702), .ZN(n_678));
   INV_X1 i_456 (.A(n_679), .ZN(n_356));
   AOI21_X1 i_457 (.A(n_19), .B1(n_18), .B2(n_714), .ZN(n_679));
   XOR2_X1 i_458 (.A(n_30), .B(n_680), .Z(n_357));
   OAI21_X1 i_459 (.A(n_733), .B1(n_736), .B2(n_731), .ZN(n_680));
   XNOR2_X1 i_460 (.A(n_687), .B(n_681), .ZN(n_358));
   NOR2_X1 i_461 (.A1(n_686), .A2(n_682), .ZN(n_681));
   INV_X1 i_462 (.A(n_683), .ZN(n_682));
   NAND3_X1 i_463 (.A1(inputB[29]), .A2(inputA[20]), .A3(n_684), .ZN(n_683));
   INV_X1 i_464 (.A(n_685), .ZN(n_684));
   NAND2_X1 i_465 (.A1(inputB[30]), .A2(inputA[21]), .ZN(n_685));
   AOI22_X1 i_466 (.A1(inputB[30]), .A2(inputA[20]), .B1(inputB[29]), .B2(
      inputA[21]), .ZN(n_686));
   AND2_X1 i_467 (.A1(inputB[31]), .A2(inputA[19]), .ZN(n_687));
   XOR2_X1 i_468 (.A(n_689), .B(n_688), .Z(n_359));
   NAND2_X1 i_469 (.A1(inputB[28]), .A2(inputA[22]), .ZN(n_688));
   OAI21_X1 i_470 (.A(n_690), .B1(n_720), .B2(n_691), .ZN(n_689));
   NAND2_X1 i_471 (.A1(n_720), .A2(n_691), .ZN(n_690));
   INV_X1 i_472 (.A(n_692), .ZN(n_691));
   NAND2_X1 i_473 (.A1(inputB[26]), .A2(inputA[24]), .ZN(n_692));
   XNOR2_X1 i_474 (.A(n_694), .B(n_693), .ZN(n_360));
   NAND2_X1 i_475 (.A1(inputB[22]), .A2(inputA[28]), .ZN(n_693));
   NOR2_X1 i_476 (.A1(n_696), .A2(n_695), .ZN(n_694));
   AOI21_X1 i_477 (.A(n_741), .B1(inputB[20]), .B2(inputA[30]), .ZN(n_695));
   INV_X1 i_478 (.A(n_697), .ZN(n_696));
   NAND3_X1 i_479 (.A1(inputB[20]), .A2(inputA[30]), .A3(n_741), .ZN(n_697));
   OAI21_X1 i_480 (.A(n_710), .B1(n_709), .B2(n_707), .ZN(n_361));
   OAI21_X1 i_481 (.A(n_728), .B1(n_730), .B2(n_726), .ZN(n_362));
   OAI21_X1 i_482 (.A(n_719), .B1(n_718), .B2(n_715), .ZN(n_363));
   OAI21_X1 i_483 (.A(n_740), .B1(n_744), .B2(n_738), .ZN(n_364));
   NAND2_X1 i_484 (.A1(inputB[19]), .A2(inputA[31]), .ZN(n_639));
   INV_X1 i_485 (.A(n_698), .ZN(n_365));
   AOI21_X1 i_486 (.A(n_11), .B1(n_10), .B2(n_699), .ZN(n_698));
   INV_X1 i_487 (.A(n_700), .ZN(n_699));
   AOI21_X1 i_488 (.A(n_5708), .B1(n_5707), .B2(n_794), .ZN(n_700));
   XOR2_X1 i_489 (.A(n_24), .B(n_701), .Z(n_366));
   XOR2_X1 i_490 (.A(n_20), .B(n_702), .Z(n_701));
   XOR2_X1 i_491 (.A(n_14), .B(n_703), .Z(n_702));
   NAND2_X1 i_492 (.A1(n_777), .A2(n_704), .ZN(n_703));
   NAND2_X1 i_493 (.A1(n_776), .A2(n_774), .ZN(n_704));
   XOR2_X1 i_494 (.A(n_22), .B(n_705), .Z(n_367));
   XOR2_X1 i_495 (.A(n_16), .B(n_706), .Z(n_705));
   XNOR2_X1 i_496 (.A(n_709), .B(n_708), .ZN(n_706));
   INV_X1 i_497 (.A(n_708), .ZN(n_707));
   AOI21_X1 i_498 (.A(n_787), .B1(n_815), .B2(n_788), .ZN(n_708));
   OAI21_X1 i_499 (.A(n_710), .B1(n_712), .B2(n_711), .ZN(n_709));
   NAND2_X1 i_500 (.A1(n_712), .A2(n_711), .ZN(n_710));
   AND2_X1 i_501 (.A1(inputB[19]), .A2(inputA[30]), .ZN(n_711));
   NAND2_X1 i_502 (.A1(inputB[18]), .A2(inputA[31]), .ZN(n_712));
   INV_X1 i_503 (.A(n_713), .ZN(n_368));
   AOI21_X1 i_504 (.A(n_7), .B1(n_6), .B2(n_751), .ZN(n_713));
   XOR2_X1 i_505 (.A(n_18), .B(n_714), .Z(n_369));
   XOR2_X1 i_506 (.A(n_716), .B(n_715), .Z(n_714));
   NAND2_X1 i_507 (.A1(inputB[28]), .A2(inputA[21]), .ZN(n_715));
   NAND2_X1 i_508 (.A1(n_719), .A2(n_717), .ZN(n_716));
   INV_X1 i_509 (.A(n_718), .ZN(n_717));
   AOI22_X1 i_510 (.A1(inputB[27]), .A2(inputA[22]), .B1(inputB[26]), .B2(
      inputA[23]), .ZN(n_718));
   NAND2_X1 i_511 (.A1(n_778), .A2(n_720), .ZN(n_719));
   INV_X1 i_512 (.A(n_721), .ZN(n_720));
   NAND2_X1 i_513 (.A1(inputB[27]), .A2(inputA[23]), .ZN(n_721));
   INV_X1 i_514 (.A(n_722), .ZN(n_370));
   AOI21_X1 i_515 (.A(n_5), .B1(n_4), .B2(n_753), .ZN(n_722));
   INV_X1 i_516 (.A(n_723), .ZN(n_371));
   AOI21_X1 i_517 (.A(n_1), .B1(n_0), .B2(n_755), .ZN(n_723));
   INV_X1 i_518 (.A(n_724), .ZN(n_372));
   AOI21_X1 i_519 (.A(n_3), .B1(n_2), .B2(n_761), .ZN(n_724));
   INV_X1 i_520 (.A(n_725), .ZN(n_373));
   AOI21_X1 i_521 (.A(n_5765), .B1(n_5764), .B2(n_772), .ZN(n_725));
   XOR2_X1 i_522 (.A(n_727), .B(n_726), .Z(n_374));
   AND2_X1 i_523 (.A1(inputB[31]), .A2(inputA[18]), .ZN(n_726));
   NAND2_X1 i_524 (.A1(n_729), .A2(n_728), .ZN(n_727));
   NAND3_X1 i_525 (.A1(inputB[30]), .A2(inputA[20]), .A3(n_767), .ZN(n_728));
   INV_X1 i_526 (.A(n_730), .ZN(n_729));
   AOI22_X1 i_527 (.A1(inputB[30]), .A2(inputA[19]), .B1(inputB[29]), .B2(
      inputA[20]), .ZN(n_730));
   XOR2_X1 i_528 (.A(n_732), .B(n_731), .Z(n_375));
   NAND2_X1 i_529 (.A1(inputB[25]), .A2(inputA[24]), .ZN(n_731));
   NAND2_X1 i_530 (.A1(n_734), .A2(n_733), .ZN(n_732));
   NAND3_X1 i_531 (.A1(inputB[24]), .A2(inputA[25]), .A3(n_737), .ZN(n_733));
   INV_X1 i_532 (.A(n_736), .ZN(n_734));
   AOI21_X1 i_533 (.A(n_737), .B1(inputB[24]), .B2(inputA[25]), .ZN(n_736));
   AND2_X1 i_534 (.A1(inputB[23]), .A2(inputA[26]), .ZN(n_737));
   XOR2_X1 i_535 (.A(n_739), .B(n_738), .Z(n_376));
   NAND2_X1 i_536 (.A1(inputB[22]), .A2(inputA[27]), .ZN(n_738));
   NAND2_X1 i_537 (.A1(n_743), .A2(n_740), .ZN(n_739));
   NAND3_X1 i_538 (.A1(inputB[20]), .A2(inputA[28]), .A3(n_741), .ZN(n_740));
   INV_X1 i_539 (.A(n_742), .ZN(n_741));
   NAND2_X1 i_540 (.A1(inputB[21]), .A2(inputA[29]), .ZN(n_742));
   INV_X1 i_541 (.A(n_744), .ZN(n_743));
   AOI22_X1 i_542 (.A1(inputB[21]), .A2(inputA[28]), .B1(inputB[20]), .B2(
      inputA[29]), .ZN(n_744));
   INV_X1 i_543 (.A(n_745), .ZN(n_5763));
   AOI21_X1 i_544 (.A(n_5760), .B1(n_5759), .B2(n_771), .ZN(n_745));
   NAND2_X1 i_545 (.A1(n_766), .A2(n_762), .ZN(n_5724));
   OAI21_X1 i_546 (.A(n_782), .B1(n_784), .B2(n_780), .ZN(n_5740));
   OAI21_X1 i_547 (.A(n_758), .B1(n_760), .B2(n_756), .ZN(n_5747));
   INV_X1 i_548 (.A(n_746), .ZN(n_5716));
   AOI21_X1 i_549 (.A(n_5713), .B1(n_5712), .B2(n_747), .ZN(n_746));
   INV_X1 i_550 (.A(n_748), .ZN(n_747));
   AOI21_X1 i_551 (.A(n_5622), .B1(n_5621), .B2(n_841), .ZN(n_748));
   XNOR2_X1 i_552 (.A(n_8), .B(n_750), .ZN(n_377));
   INV_X1 i_553 (.A(n_750), .ZN(n_749));
   AOI21_X1 i_554 (.A(n_5703), .B1(n_5702), .B2(n_797), .ZN(n_750));
   XNOR2_X1 i_555 (.A(n_6), .B(n_752), .ZN(n_378));
   INV_X1 i_556 (.A(n_752), .ZN(n_751));
   AOI21_X1 i_557 (.A(n_5693), .B1(n_5692), .B2(n_800), .ZN(n_752));
   XNOR2_X1 i_558 (.A(n_4), .B(n_754), .ZN(n_379));
   INV_X1 i_559 (.A(n_754), .ZN(n_753));
   AOI21_X1 i_560 (.A(n_5688), .B1(n_5687), .B2(n_802), .ZN(n_754));
   XOR2_X1 i_561 (.A(n_0), .B(n_755), .Z(n_380));
   XOR2_X1 i_562 (.A(n_757), .B(n_756), .Z(n_755));
   NAND2_X1 i_563 (.A1(inputB[22]), .A2(inputA[26]), .ZN(n_756));
   NAND2_X1 i_564 (.A1(n_759), .A2(n_758), .ZN(n_757));
   NAND3_X1 i_565 (.A1(inputB[21]), .A2(inputA[28]), .A3(n_835), .ZN(n_758));
   INV_X1 i_566 (.A(n_760), .ZN(n_759));
   AOI22_X1 i_567 (.A1(inputB[21]), .A2(inputA[27]), .B1(inputB[20]), .B2(
      inputA[28]), .ZN(n_760));
   XOR2_X1 i_568 (.A(n_2), .B(n_761), .Z(n_381));
   XNOR2_X1 i_569 (.A(n_764), .B(n_763), .ZN(n_761));
   NAND2_X1 i_570 (.A1(n_765), .A2(n_763), .ZN(n_762));
   NAND2_X1 i_571 (.A1(inputB[31]), .A2(inputA[17]), .ZN(n_763));
   NAND2_X1 i_572 (.A1(n_766), .A2(n_765), .ZN(n_764));
   NAND2_X1 i_573 (.A1(n_825), .A2(n_768), .ZN(n_765));
   NAND2_X1 i_574 (.A1(n_824), .A2(n_767), .ZN(n_766));
   INV_X1 i_575 (.A(n_768), .ZN(n_767));
   NAND2_X1 i_576 (.A1(inputB[29]), .A2(inputA[19]), .ZN(n_768));
   INV_X1 i_577 (.A(n_769), .ZN(n_5701));
   AOI21_X1 i_578 (.A(n_5698), .B1(n_5697), .B2(n_795), .ZN(n_769));
   INV_X1 i_579 (.A(n_770), .ZN(n_5686));
   AOI21_X1 i_580 (.A(n_5683), .B1(n_5682), .B2(n_811), .ZN(n_770));
   XOR2_X1 i_581 (.A(n_5759), .B(n_771), .Z(n_5761));
   OAI21_X1 i_582 (.A(n_828), .B1(n_830), .B2(n_826), .ZN(n_771));
   XNOR2_X1 i_583 (.A(n_5764), .B(n_773), .ZN(n_5766));
   INV_X1 i_584 (.A(n_773), .ZN(n_772));
   AOI21_X1 i_585 (.A(n_5678), .B1(n_5677), .B2(n_801), .ZN(n_773));
   XOR2_X1 i_586 (.A(n_775), .B(n_774), .Z(n_5732));
   AND2_X1 i_587 (.A1(inputB[28]), .A2(inputA[20]), .ZN(n_774));
   AND2_X1 i_588 (.A1(n_777), .A2(n_776), .ZN(n_775));
   NAND2_X1 i_589 (.A1(n_807), .A2(n_779), .ZN(n_776));
   NAND2_X1 i_590 (.A1(n_806), .A2(n_778), .ZN(n_777));
   INV_X1 i_591 (.A(n_779), .ZN(n_778));
   NAND2_X1 i_592 (.A1(inputB[26]), .A2(inputA[22]), .ZN(n_779));
   XOR2_X1 i_593 (.A(n_781), .B(n_780), .Z(n_5739));
   NAND2_X1 i_594 (.A1(inputB[25]), .A2(inputA[23]), .ZN(n_780));
   NAND2_X1 i_595 (.A1(n_783), .A2(n_782), .ZN(n_781));
   NAND4_X1 i_596 (.A1(inputB[24]), .A2(inputA[24]), .A3(inputB[23]), .A4(
      inputA[25]), .ZN(n_782));
   INV_X1 i_597 (.A(n_784), .ZN(n_783));
   AOI22_X1 i_598 (.A1(inputB[24]), .A2(inputA[24]), .B1(inputB[23]), .B2(
      inputA[25]), .ZN(n_784));
   XOR2_X1 i_599 (.A(n_815), .B(n_785), .Z(n_5752));
   NAND2_X1 i_600 (.A1(n_788), .A2(n_786), .ZN(n_785));
   INV_X1 i_601 (.A(n_787), .ZN(n_786));
   AOI211_X1 i_602 (.A(n_5762), .B(n_5753), .C1(inputB[19]), .C2(inputA[29]), 
      .ZN(n_787));
   OAI211_X1 i_603 (.A(inputB[19]), .B(inputA[29]), .C1(n_5762), .C2(n_5753), 
      .ZN(n_788));
   INV_X1 i_604 (.A(n_789), .ZN(n_5676));
   AOI21_X1 i_605 (.A(n_5673), .B1(n_5672), .B2(n_819), .ZN(n_789));
   NOR2_X1 i_606 (.A1(n_823), .A2(n_790), .ZN(n_5638));
   AOI21_X1 i_607 (.A(n_821), .B1(n_872), .B2(n_824), .ZN(n_790));
   OAI21_X1 i_608 (.A(n_805), .B1(n_809), .B2(n_808), .ZN(n_5647));
   AOI22_X1 i_609 (.A1(n_883), .A2(n_836), .B1(n_834), .B2(n_832), .ZN(n_5661));
   OAI21_X1 i_610 (.A(n_814), .B1(n_816), .B2(n_812), .ZN(n_5668));
   INV_X1 i_611 (.A(n_791), .ZN(n_5630));
   AOI21_X1 i_612 (.A(n_5627), .B1(n_5626), .B2(n_792), .ZN(n_791));
   INV_X1 i_613 (.A(n_793), .ZN(n_792));
   AOI21_X1 i_614 (.A(n_5528), .B1(n_5527), .B2(n_898), .ZN(n_793));
   XOR2_X1 i_615 (.A(n_5707), .B(n_794), .Z(n_5709));
   XNOR2_X1 i_616 (.A(n_5697), .B(n_796), .ZN(n_794));
   INV_X1 i_617 (.A(n_796), .ZN(n_795));
   AOI21_X1 i_618 (.A(n_5597), .B1(n_5596), .B2(n_845), .ZN(n_796));
   XNOR2_X1 i_619 (.A(n_5702), .B(n_798), .ZN(n_5704));
   INV_X1 i_620 (.A(n_798), .ZN(n_797));
   AOI21_X1 i_621 (.A(n_5612), .B1(n_5611), .B2(n_853), .ZN(n_798));
   INV_X1 i_622 (.A(n_799), .ZN(n_5620));
   AOI21_X1 i_623 (.A(n_5617), .B1(n_5616), .B2(n_844), .ZN(n_799));
   XOR2_X1 i_624 (.A(n_5692), .B(n_800), .Z(n_5694));
   XOR2_X1 i_625 (.A(n_5677), .B(n_801), .Z(n_800));
   NAND2_X1 i_626 (.A1(n_871), .A2(n_867), .ZN(n_801));
   XOR2_X1 i_627 (.A(n_5687), .B(n_802), .Z(n_5689));
   XNOR2_X1 i_628 (.A(n_809), .B(n_803), .ZN(n_802));
   NOR2_X1 i_629 (.A1(n_808), .A2(n_804), .ZN(n_803));
   INV_X1 i_630 (.A(n_805), .ZN(n_804));
   NAND3_X1 i_631 (.A1(inputB[26]), .A2(inputA[20]), .A3(n_806), .ZN(n_805));
   INV_X1 i_632 (.A(n_807), .ZN(n_806));
   NAND2_X1 i_633 (.A1(inputB[27]), .A2(inputA[21]), .ZN(n_807));
   AOI22_X1 i_634 (.A1(inputB[27]), .A2(inputA[20]), .B1(inputB[26]), .B2(
      inputA[21]), .ZN(n_808));
   NAND2_X1 i_635 (.A1(inputB[28]), .A2(inputA[19]), .ZN(n_809));
   INV_X1 i_636 (.A(n_810), .ZN(n_5610));
   AOI21_X1 i_637 (.A(n_5607), .B1(n_5606), .B2(n_842), .ZN(n_810));
   XOR2_X1 i_638 (.A(n_5682), .B(n_811), .Z(n_5684));
   XOR2_X1 i_639 (.A(n_813), .B(n_812), .Z(n_811));
   NAND2_X1 i_640 (.A1(inputB[19]), .A2(inputA[28]), .ZN(n_812));
   NAND2_X1 i_641 (.A1(n_817), .A2(n_814), .ZN(n_813));
   OR3_X1 i_642 (.A1(n_5762), .A2(n_5750), .A3(n_815), .ZN(n_814));
   NAND2_X1 i_643 (.A1(inputB[18]), .A2(inputA[30]), .ZN(n_815));
   INV_X1 i_644 (.A(n_817), .ZN(n_816));
   OAI21_X1 i_645 (.A(n_851), .B1(n_5762), .B2(n_5751), .ZN(n_817));
   INV_X1 i_646 (.A(n_818), .ZN(n_5605));
   AOI21_X1 i_647 (.A(n_5602), .B1(n_5601), .B2(n_856), .ZN(n_818));
   XOR2_X1 i_648 (.A(n_5672), .B(n_819), .Z(n_5674));
   OAI21_X1 i_649 (.A(n_881), .B1(n_885), .B2(n_879), .ZN(n_819));
   INV_X1 i_650 (.A(n_820), .ZN(n_5595));
   AOI21_X1 i_651 (.A(n_5592), .B1(n_5591), .B2(n_865), .ZN(n_820));
   XOR2_X1 i_652 (.A(n_822), .B(n_821), .Z(n_5637));
   NAND2_X1 i_653 (.A1(inputB[31]), .A2(inputA[16]), .ZN(n_821));
   AOI21_X1 i_654 (.A(n_823), .B1(n_872), .B2(n_824), .ZN(n_822));
   AOI22_X1 i_655 (.A1(inputB[30]), .A2(inputA[17]), .B1(inputB[29]), .B2(
      inputA[18]), .ZN(n_823));
   INV_X1 i_656 (.A(n_825), .ZN(n_824));
   NAND2_X1 i_657 (.A1(inputB[30]), .A2(inputA[18]), .ZN(n_825));
   XOR2_X1 i_658 (.A(n_827), .B(n_826), .Z(n_5653));
   NAND2_X1 i_659 (.A1(inputB[25]), .A2(inputA[22]), .ZN(n_826));
   NAND2_X1 i_660 (.A1(n_829), .A2(n_828), .ZN(n_827));
   NAND4_X1 i_661 (.A1(inputB[24]), .A2(inputA[23]), .A3(inputB[23]), .A4(
      inputA[24]), .ZN(n_828));
   INV_X1 i_662 (.A(n_830), .ZN(n_829));
   AOI22_X1 i_663 (.A1(inputB[24]), .A2(inputA[23]), .B1(inputB[23]), .B2(
      inputA[24]), .ZN(n_830));
   XOR2_X1 i_664 (.A(n_833), .B(n_832), .Z(n_5660));
   NAND2_X1 i_665 (.A1(inputB[22]), .A2(inputA[25]), .ZN(n_832));
   OAI21_X1 i_666 (.A(n_834), .B1(n_882), .B2(n_835), .ZN(n_833));
   NAND2_X1 i_667 (.A1(n_882), .A2(n_835), .ZN(n_834));
   INV_X1 i_668 (.A(n_836), .ZN(n_835));
   NAND2_X1 i_669 (.A1(inputB[20]), .A2(inputA[27]), .ZN(n_836));
   AOI21_X1 i_670 (.A(n_888), .B1(n_889), .B2(n_886), .ZN(n_5581));
   INV_X1 i_671 (.A(n_837), .ZN(n_5590));
   AOI21_X1 i_672 (.A(n_5587), .B1(n_5586), .B2(n_843), .ZN(n_837));
   OAI21_X1 i_673 (.A(n_859), .B1(n_861), .B2(n_857), .ZN(n_5553));
   OAI21_X1 i_674 (.A(n_876), .B1(n_878), .B2(n_874), .ZN(n_5560));
   OAI21_X1 i_675 (.A(n_850), .B1(n_849), .B2(n_846), .ZN(n_5574));
   NAND2_X1 i_676 (.A1(inputB[16]), .A2(inputA[31]), .ZN(n_543));
   INV_X1 i_677 (.A(n_838), .ZN(n_5536));
   AOI21_X1 i_678 (.A(n_5533), .B1(n_5532), .B2(n_839), .ZN(n_838));
   INV_X1 i_679 (.A(n_840), .ZN(n_839));
   AOI21_X1 i_680 (.A(n_5429), .B1(n_5428), .B2(n_955), .ZN(n_840));
   XOR2_X1 i_681 (.A(n_5621), .B(n_841), .Z(n_5623));
   XOR2_X1 i_682 (.A(n_5606), .B(n_842), .Z(n_841));
   XOR2_X1 i_683 (.A(n_5586), .B(n_843), .Z(n_842));
   AOI21_X1 i_684 (.A(n_906), .B1(n_907), .B2(n_903), .ZN(n_843));
   XOR2_X1 i_685 (.A(n_5616), .B(n_844), .Z(n_5618));
   XOR2_X1 i_686 (.A(n_5596), .B(n_845), .Z(n_844));
   XOR2_X1 i_687 (.A(n_847), .B(n_846), .Z(n_845));
   NAND2_X1 i_688 (.A1(inputB[19]), .A2(inputA[27]), .ZN(n_846));
   NAND2_X1 i_689 (.A1(n_850), .A2(n_848), .ZN(n_847));
   INV_X1 i_690 (.A(n_849), .ZN(n_848));
   AOI22_X1 i_691 (.A1(inputB[18]), .A2(inputA[28]), .B1(inputB[17]), .B2(
      inputA[29]), .ZN(n_849));
   OR2_X1 i_692 (.A1(n_949), .A2(n_851), .ZN(n_850));
   NAND2_X1 i_693 (.A1(inputB[18]), .A2(inputA[29]), .ZN(n_851));
   INV_X1 i_694 (.A(n_852), .ZN(n_5526));
   AOI21_X1 i_695 (.A(n_5523), .B1(n_5522), .B2(n_901), .ZN(n_852));
   XNOR2_X1 i_696 (.A(n_5611), .B(n_854), .ZN(n_5613));
   INV_X1 i_697 (.A(n_854), .ZN(n_853));
   AOI21_X1 i_698 (.A(n_5508), .B1(n_5507), .B2(n_913), .ZN(n_854));
   INV_X1 i_699 (.A(n_855), .ZN(n_5521));
   AOI21_X1 i_700 (.A(n_5518), .B1(n_5517), .B2(n_899), .ZN(n_855));
   XOR2_X1 i_701 (.A(n_5601), .B(n_856), .Z(n_5603));
   XOR2_X1 i_702 (.A(n_858), .B(n_857), .Z(n_856));
   NAND2_X1 i_703 (.A1(inputB[28]), .A2(inputA[18]), .ZN(n_857));
   NAND2_X1 i_704 (.A1(n_860), .A2(n_859), .ZN(n_858));
   NAND3_X1 i_705 (.A1(inputB[27]), .A2(inputA[20]), .A3(n_937), .ZN(n_859));
   INV_X1 i_706 (.A(n_861), .ZN(n_860));
   AOI22_X1 i_707 (.A1(inputB[27]), .A2(inputA[19]), .B1(inputB[26]), .B2(
      inputA[20]), .ZN(n_861));
   INV_X1 i_708 (.A(n_862), .ZN(n_5516));
   AOI21_X1 i_709 (.A(n_5513), .B1(n_5512), .B2(n_911), .ZN(n_862));
   INV_X1 i_710 (.A(n_863), .ZN(n_5501));
   AOI21_X1 i_711 (.A(n_5498), .B1(n_5497), .B2(n_916), .ZN(n_863));
   INV_X1 i_712 (.A(n_864), .ZN(n_5506));
   AOI21_X1 i_713 (.A(n_5503), .B1(n_5502), .B2(n_902), .ZN(n_864));
   XNOR2_X1 i_714 (.A(n_5591), .B(n_866), .ZN(n_5593));
   INV_X1 i_715 (.A(n_866), .ZN(n_865));
   AOI21_X1 i_716 (.A(n_5493), .B1(n_5492), .B2(n_925), .ZN(n_866));
   XNOR2_X1 i_717 (.A(n_869), .B(n_868), .ZN(n_5543));
   NAND2_X1 i_718 (.A1(n_870), .A2(n_868), .ZN(n_867));
   NAND2_X1 i_719 (.A1(inputB[31]), .A2(inputA[15]), .ZN(n_868));
   NAND2_X1 i_720 (.A1(n_871), .A2(n_870), .ZN(n_869));
   NAND2_X1 i_721 (.A1(n_932), .A2(n_873), .ZN(n_870));
   NAND2_X1 i_722 (.A1(n_931), .A2(n_872), .ZN(n_871));
   INV_X1 i_723 (.A(n_873), .ZN(n_872));
   NAND2_X1 i_724 (.A1(inputB[29]), .A2(inputA[17]), .ZN(n_873));
   XOR2_X1 i_725 (.A(n_875), .B(n_874), .Z(n_5559));
   NAND2_X1 i_726 (.A1(inputB[25]), .A2(inputA[21]), .ZN(n_874));
   NAND2_X1 i_727 (.A1(n_877), .A2(n_876), .ZN(n_875));
   NAND3_X1 i_728 (.A1(inputB[23]), .A2(inputA[23]), .A3(n_908), .ZN(n_876));
   INV_X1 i_729 (.A(n_878), .ZN(n_877));
   AOI21_X1 i_730 (.A(n_908), .B1(inputB[23]), .B2(inputA[23]), .ZN(n_878));
   XOR2_X1 i_731 (.A(n_880), .B(n_879), .Z(n_5566));
   NAND2_X1 i_732 (.A1(inputB[22]), .A2(inputA[24]), .ZN(n_879));
   NAND2_X1 i_733 (.A1(n_884), .A2(n_881), .ZN(n_880));
   NAND2_X1 i_734 (.A1(n_944), .A2(n_882), .ZN(n_881));
   INV_X1 i_735 (.A(n_883), .ZN(n_882));
   NAND2_X1 i_736 (.A1(inputB[21]), .A2(inputA[26]), .ZN(n_883));
   INV_X1 i_737 (.A(n_885), .ZN(n_884));
   AOI22_X1 i_738 (.A1(inputB[21]), .A2(inputA[25]), .B1(inputB[20]), .B2(
      inputA[26]), .ZN(n_885));
   XNOR2_X1 i_739 (.A(n_887), .B(n_886), .ZN(n_5580));
   AOI21_X1 i_740 (.A(n_921), .B1(n_919), .B2(n_917), .ZN(n_886));
   NOR2_X1 i_741 (.A1(n_890), .A2(n_888), .ZN(n_887));
   AND3_X1 i_742 (.A1(inputB[15]), .A2(inputA[31]), .A3(n_922), .ZN(n_888));
   INV_X1 i_743 (.A(n_890), .ZN(n_889));
   AOI21_X1 i_744 (.A(n_922), .B1(inputB[15]), .B2(inputA[31]), .ZN(n_890));
   INV_X1 i_745 (.A(n_891), .ZN(n_5491));
   AOI21_X1 i_746 (.A(n_5488), .B1(n_5487), .B2(n_924), .ZN(n_891));
   INV_X1 i_747 (.A(n_892), .ZN(n_5445));
   AOI22_X1 i_748 (.A1(n_993), .A2(n_931), .B1(n_929), .B2(n_928), .ZN(n_892));
   NAND2_X1 i_749 (.A1(n_936), .A2(n_893), .ZN(n_5454));
   NAND2_X1 i_750 (.A1(n_935), .A2(n_933), .ZN(n_893));
   OAI21_X1 i_751 (.A(n_941), .B1(n_943), .B2(n_939), .ZN(n_5468));
   NAND2_X1 i_752 (.A1(n_948), .A2(n_894), .ZN(n_5475));
   NAND2_X1 i_753 (.A1(n_947), .A2(n_945), .ZN(n_894));
   INV_X1 i_754 (.A(n_895), .ZN(n_5437));
   AOI21_X1 i_755 (.A(n_5434), .B1(n_5433), .B2(n_896), .ZN(n_895));
   INV_X1 i_756 (.A(n_897), .ZN(n_896));
   AOI21_X1 i_757 (.A(n_5326), .B1(n_5325), .B2(n_1015), .ZN(n_897));
   XOR2_X1 i_758 (.A(n_5527), .B(n_898), .Z(n_5529));
   XNOR2_X1 i_759 (.A(n_5517), .B(n_900), .ZN(n_898));
   INV_X1 i_760 (.A(n_900), .ZN(n_899));
   AOI21_X1 i_761 (.A(n_5414), .B1(n_5413), .B2(n_966), .ZN(n_900));
   XOR2_X1 i_762 (.A(n_5522), .B(n_901), .Z(n_5524));
   XOR2_X1 i_763 (.A(n_5502), .B(n_902), .Z(n_901));
   XOR2_X1 i_764 (.A(n_904), .B(n_903), .Z(n_902));
   NAND2_X1 i_765 (.A1(inputB[25]), .A2(inputA[20]), .ZN(n_903));
   NAND2_X1 i_766 (.A1(n_907), .A2(n_905), .ZN(n_904));
   INV_X1 i_767 (.A(n_906), .ZN(n_905));
   AOI22_X1 i_768 (.A1(inputB[24]), .A2(inputA[21]), .B1(inputB[23]), .B2(
      inputA[22]), .ZN(n_906));
   NAND2_X1 i_769 (.A1(n_998), .A2(n_908), .ZN(n_907));
   AND2_X1 i_770 (.A1(inputB[24]), .A2(inputA[22]), .ZN(n_908));
   INV_X1 i_771 (.A(n_909), .ZN(n_5427));
   AOI21_X1 i_772 (.A(n_5424), .B1(n_5423), .B2(n_965), .ZN(n_909));
   INV_X1 i_773 (.A(n_910), .ZN(n_5422));
   AOI21_X1 i_774 (.A(n_5419), .B1(n_5418), .B2(n_956), .ZN(n_910));
   XNOR2_X1 i_775 (.A(n_5512), .B(n_912), .ZN(n_5514));
   INV_X1 i_776 (.A(n_912), .ZN(n_911));
   AOI21_X1 i_777 (.A(n_5404), .B1(n_5403), .B2(n_957), .ZN(n_912));
   XNOR2_X1 i_778 (.A(n_5507), .B(n_914), .ZN(n_5509));
   INV_X1 i_779 (.A(n_914), .ZN(n_913));
   AOI21_X1 i_780 (.A(n_5394), .B1(n_5393), .B2(n_982), .ZN(n_914));
   INV_X1 i_781 (.A(n_915), .ZN(n_5412));
   AOI21_X1 i_782 (.A(n_5409), .B1(n_5408), .B2(n_970), .ZN(n_915));
   XOR2_X1 i_783 (.A(n_5497), .B(n_916), .Z(n_5499));
   XOR2_X1 i_784 (.A(n_918), .B(n_917), .Z(n_916));
   NAND2_X1 i_785 (.A1(inputB[14]), .A2(inputA[31]), .ZN(n_917));
   NOR2_X1 i_786 (.A1(n_921), .A2(n_920), .ZN(n_918));
   INV_X1 i_787 (.A(n_920), .ZN(n_919));
   AOI22_X1 i_788 (.A1(inputB[15]), .A2(inputA[30]), .B1(inputB[16]), .B2(
      inputA[29]), .ZN(n_920));
   NOR2_X1 i_789 (.A1(n_1100), .A2(n_922), .ZN(n_921));
   NAND2_X1 i_790 (.A1(inputB[16]), .A2(inputA[30]), .ZN(n_922));
   INV_X1 i_791 (.A(n_923), .ZN(n_5402));
   AOI21_X1 i_792 (.A(n_5399), .B1(n_5398), .B2(n_974), .ZN(n_923));
   XOR2_X1 i_793 (.A(n_5487), .B(n_924), .Z(n_5489));
   OAI21_X1 i_794 (.A(n_1002), .B1(n_1004), .B2(n_1000), .ZN(n_924));
   XOR2_X1 i_795 (.A(n_5492), .B(n_925), .Z(n_5494));
   NAND2_X1 i_796 (.A1(n_992), .A2(n_926), .ZN(n_925));
   NAND2_X1 i_797 (.A1(n_990), .A2(n_988), .ZN(n_926));
   XOR2_X1 i_798 (.A(n_929), .B(n_928), .Z(n_5444));
   NAND2_X1 i_799 (.A1(inputB[31]), .A2(inputA[14]), .ZN(n_928));
   AOI21_X1 i_800 (.A(n_930), .B1(n_993), .B2(n_931), .ZN(n_929));
   AOI22_X1 i_801 (.A1(inputB[30]), .A2(inputA[15]), .B1(inputB[29]), .B2(
      inputA[16]), .ZN(n_930));
   INV_X1 i_802 (.A(n_932), .ZN(n_931));
   NAND2_X1 i_803 (.A1(inputB[30]), .A2(inputA[16]), .ZN(n_932));
   XOR2_X1 i_804 (.A(n_934), .B(n_933), .Z(n_5453));
   AND2_X1 i_805 (.A1(inputB[28]), .A2(inputA[17]), .ZN(n_933));
   AND2_X1 i_806 (.A1(n_936), .A2(n_935), .ZN(n_934));
   NAND2_X1 i_807 (.A1(n_964), .A2(n_938), .ZN(n_935));
   NAND2_X1 i_808 (.A1(n_963), .A2(n_937), .ZN(n_936));
   INV_X1 i_809 (.A(n_938), .ZN(n_937));
   NAND2_X1 i_810 (.A1(inputB[26]), .A2(inputA[19]), .ZN(n_938));
   XOR2_X1 i_811 (.A(n_940), .B(n_939), .Z(n_5467));
   NAND2_X1 i_812 (.A1(inputB[22]), .A2(inputA[23]), .ZN(n_939));
   NAND2_X1 i_813 (.A1(n_942), .A2(n_941), .ZN(n_940));
   NAND3_X1 i_814 (.A1(inputB[21]), .A2(inputA[24]), .A3(n_944), .ZN(n_941));
   INV_X1 i_815 (.A(n_943), .ZN(n_942));
   AOI21_X1 i_816 (.A(n_944), .B1(inputB[21]), .B2(inputA[24]), .ZN(n_943));
   AND2_X1 i_817 (.A1(inputB[20]), .A2(inputA[25]), .ZN(n_944));
   XOR2_X1 i_818 (.A(n_946), .B(n_945), .Z(n_5474));
   AND2_X1 i_819 (.A1(inputB[19]), .A2(inputA[26]), .ZN(n_945));
   AND2_X1 i_820 (.A1(n_948), .A2(n_947), .ZN(n_946));
   NAND2_X1 i_821 (.A1(n_980), .A2(n_949), .ZN(n_947));
   OR2_X1 i_822 (.A1(n_980), .A2(n_949), .ZN(n_948));
   NAND2_X1 i_823 (.A1(inputB[17]), .A2(inputA[28]), .ZN(n_949));
   INV_X1 i_824 (.A(n_950), .ZN(n_5387));
   AOI21_X1 i_825 (.A(n_5384), .B1(n_5383), .B2(n_971), .ZN(n_950));
   INV_X1 i_826 (.A(n_951), .ZN(n_5392));
   AOI21_X1 i_827 (.A(n_5389), .B1(n_5388), .B2(n_986), .ZN(n_951));
   OAI21_X1 i_828 (.A(n_962), .B1(n_961), .B2(n_958), .ZN(n_5351));
   AOI22_X1 i_829 (.A1(n_1081), .A2(n_999), .B1(n_997), .B2(n_995), .ZN(n_5358));
   OAI21_X1 i_830 (.A(n_979), .B1(n_978), .B2(n_975), .ZN(n_5372));
   OAI21_X1 i_831 (.A(n_1009), .B1(n_1007), .B2(n_1005), .ZN(n_5379));
   INV_X1 i_832 (.A(n_952), .ZN(n_5334));
   AOI21_X1 i_833 (.A(n_5331), .B1(n_5330), .B2(n_953), .ZN(n_952));
   INV_X1 i_834 (.A(n_954), .ZN(n_953));
   AOI21_X1 i_835 (.A(n_5215), .B1(n_5214), .B2(n_1110), .ZN(n_954));
   XOR2_X1 i_836 (.A(n_5428), .B(n_955), .Z(n_5430));
   XOR2_X1 i_837 (.A(n_5418), .B(n_956), .Z(n_955));
   XOR2_X1 i_838 (.A(n_5403), .B(n_957), .Z(n_956));
   XOR2_X1 i_839 (.A(n_959), .B(n_958), .Z(n_957));
   NAND2_X1 i_840 (.A1(inputB[28]), .A2(inputA[16]), .ZN(n_958));
   NAND2_X1 i_841 (.A1(n_962), .A2(n_960), .ZN(n_959));
   INV_X1 i_842 (.A(n_961), .ZN(n_960));
   AOI22_X1 i_843 (.A1(inputB[27]), .A2(inputA[17]), .B1(inputB[26]), .B2(
      inputA[18]), .ZN(n_961));
   NAND2_X1 i_844 (.A1(n_1067), .A2(n_963), .ZN(n_962));
   INV_X1 i_845 (.A(n_964), .ZN(n_963));
   NAND2_X1 i_846 (.A1(inputB[27]), .A2(inputA[18]), .ZN(n_964));
   XOR2_X1 i_847 (.A(n_5423), .B(n_965), .Z(n_5425));
   XNOR2_X1 i_848 (.A(n_5413), .B(n_967), .ZN(n_965));
   INV_X1 i_849 (.A(n_967), .ZN(n_966));
   AOI21_X1 i_850 (.A(n_5291), .B1(n_5290), .B2(n_1026), .ZN(n_967));
   INV_X1 i_851 (.A(n_968), .ZN(n_5324));
   AOI21_X1 i_852 (.A(n_5321), .B1(n_5320), .B2(n_1024), .ZN(n_968));
   INV_X1 i_853 (.A(n_969), .ZN(n_5319));
   AOI21_X1 i_854 (.A(n_5316), .B1(n_5315), .B2(n_1016), .ZN(n_969));
   XOR2_X1 i_855 (.A(n_5408), .B(n_970), .Z(n_5410));
   XOR2_X1 i_856 (.A(n_5383), .B(n_971), .Z(n_970));
   NAND2_X1 i_857 (.A1(n_1088), .A2(n_972), .ZN(n_971));
   NAND2_X1 i_858 (.A1(n_1087), .A2(n_1085), .ZN(n_972));
   INV_X1 i_859 (.A(n_973), .ZN(n_5314));
   AOI21_X1 i_860 (.A(n_5311), .B1(n_5310), .B2(n_1025), .ZN(n_973));
   XOR2_X1 i_861 (.A(n_5398), .B(n_974), .Z(n_5400));
   XOR2_X1 i_862 (.A(n_976), .B(n_975), .Z(n_974));
   NAND2_X1 i_863 (.A1(inputB[19]), .A2(inputA[25]), .ZN(n_975));
   NAND2_X1 i_864 (.A1(n_979), .A2(n_977), .ZN(n_976));
   INV_X1 i_865 (.A(n_978), .ZN(n_977));
   AOI22_X1 i_866 (.A1(inputB[18]), .A2(inputA[26]), .B1(inputB[17]), .B2(
      inputA[27]), .ZN(n_978));
   OR2_X1 i_867 (.A1(n_1089), .A2(n_980), .ZN(n_979));
   NAND2_X1 i_868 (.A1(inputB[18]), .A2(inputA[27]), .ZN(n_980));
   INV_X1 i_869 (.A(n_981), .ZN(n_5309));
   AOI21_X1 i_870 (.A(n_5306), .B1(n_5305), .B2(n_1038), .ZN(n_981));
   XNOR2_X1 i_871 (.A(n_5393), .B(n_983), .ZN(n_5395));
   INV_X1 i_872 (.A(n_983), .ZN(n_982));
   AOI21_X1 i_873 (.A(n_5281), .B1(n_5280), .B2(n_1041), .ZN(n_983));
   INV_X1 i_874 (.A(n_984), .ZN(n_5299));
   AOI21_X1 i_875 (.A(n_5296), .B1(n_5295), .B2(n_1044), .ZN(n_984));
   INV_X1 i_876 (.A(n_985), .ZN(n_5304));
   AOI21_X1 i_877 (.A(n_5301), .B1(n_5300), .B2(n_1017), .ZN(n_985));
   XOR2_X1 i_878 (.A(n_5388), .B(n_986), .Z(n_5390));
   NAND2_X1 i_879 (.A1(n_1066), .A2(n_987), .ZN(n_986));
   NAND2_X1 i_880 (.A1(n_1065), .A2(n_1063), .ZN(n_987));
   XOR2_X1 i_881 (.A(n_989), .B(n_988), .Z(n_5341));
   NAND2_X1 i_882 (.A1(inputB[31]), .A2(inputA[13]), .ZN(n_988));
   AND2_X1 i_883 (.A1(n_992), .A2(n_990), .ZN(n_989));
   NAND2_X1 i_884 (.A1(n_1023), .A2(n_994), .ZN(n_990));
   NAND2_X1 i_885 (.A1(n_1021), .A2(n_993), .ZN(n_992));
   INV_X1 i_886 (.A(n_994), .ZN(n_993));
   NAND2_X1 i_887 (.A1(inputB[29]), .A2(inputA[15]), .ZN(n_994));
   XOR2_X1 i_888 (.A(n_996), .B(n_995), .Z(n_5357));
   NAND2_X1 i_889 (.A1(inputB[25]), .A2(inputA[19]), .ZN(n_995));
   OAI21_X1 i_890 (.A(n_997), .B1(n_1080), .B2(n_998), .ZN(n_996));
   NAND2_X1 i_891 (.A1(n_1080), .A2(n_998), .ZN(n_997));
   INV_X1 i_892 (.A(n_999), .ZN(n_998));
   NAND2_X1 i_893 (.A1(inputB[23]), .A2(inputA[21]), .ZN(n_999));
   XOR2_X1 i_894 (.A(n_1001), .B(n_1000), .Z(n_5364));
   NAND2_X1 i_895 (.A1(inputB[22]), .A2(inputA[22]), .ZN(n_1000));
   NAND2_X1 i_896 (.A1(n_1003), .A2(n_1002), .ZN(n_1001));
   NAND3_X1 i_897 (.A1(inputB[20]), .A2(inputA[24]), .A3(n_1054), .ZN(n_1002));
   INV_X1 i_898 (.A(n_1004), .ZN(n_1003));
   AOI21_X1 i_899 (.A(n_1054), .B1(inputB[20]), .B2(inputA[24]), .ZN(n_1004));
   XNOR2_X1 i_900 (.A(n_1006), .B(n_1005), .ZN(n_5378));
   NAND2_X1 i_901 (.A1(inputB[16]), .A2(inputA[28]), .ZN(n_1005));
   NOR2_X1 i_902 (.A1(n_1008), .A2(n_1007), .ZN(n_1006));
   AOI21_X1 i_903 (.A(n_1096), .B1(inputB[14]), .B2(inputA[30]), .ZN(n_1007));
   INV_X1 i_904 (.A(n_1009), .ZN(n_1008));
   NAND3_X1 i_905 (.A1(inputB[14]), .A2(inputA[30]), .A3(n_1096), .ZN(n_1009));
   OAI21_X1 i_906 (.A(n_1032), .B1(n_1031), .B2(n_1027), .ZN(n_5275));
   INV_X1 i_907 (.A(n_1010), .ZN(n_5289));
   AOI21_X1 i_908 (.A(n_5286), .B1(n_5285), .B2(n_1060), .ZN(n_1010));
   INV_X1 i_909 (.A(n_1011), .ZN(n_5231));
   AOI22_X1 i_910 (.A1(n_1181), .A2(n_1021), .B1(n_1019), .B2(n_1018), .ZN(
      n_1011));
   OAI21_X1 i_911 (.A(n_1079), .B1(n_1083), .B2(n_1075), .ZN(n_5247));
   OAI21_X1 i_912 (.A(n_1051), .B1(n_1050), .B2(n_1047), .ZN(n_5254));
   OAI21_X1 i_913 (.A(n_1095), .B1(n_1094), .B2(n_1090), .ZN(n_5268));
   NAND2_X1 i_914 (.A1(inputB[13]), .A2(inputA[31]), .ZN(n_447));
   INV_X1 i_915 (.A(n_1012), .ZN(n_5223));
   AOI21_X1 i_916 (.A(n_5220), .B1(n_5219), .B2(n_1013), .ZN(n_1012));
   INV_X1 i_917 (.A(n_1014), .ZN(n_1013));
   AOI21_X1 i_918 (.A(n_5099), .B1(n_5098), .B2(n_1222), .ZN(n_1014));
   XOR2_X1 i_919 (.A(n_5325), .B(n_1015), .Z(n_5327));
   XOR2_X1 i_920 (.A(n_5315), .B(n_1016), .Z(n_1015));
   XOR2_X1 i_921 (.A(n_5300), .B(n_1017), .Z(n_1016));
   XOR2_X1 i_922 (.A(n_1019), .B(n_1018), .Z(n_1017));
   NAND2_X1 i_923 (.A1(inputB[31]), .A2(inputA[12]), .ZN(n_1018));
   AOI21_X1 i_924 (.A(n_1020), .B1(n_1181), .B2(n_1021), .ZN(n_1019));
   AOI22_X1 i_925 (.A1(inputB[30]), .A2(inputA[13]), .B1(inputB[29]), .B2(
      inputA[14]), .ZN(n_1020));
   INV_X1 i_926 (.A(n_1023), .ZN(n_1021));
   NAND2_X1 i_927 (.A1(inputB[30]), .A2(inputA[14]), .ZN(n_1023));
   XOR2_X1 i_928 (.A(n_5320), .B(n_1024), .Z(n_5322));
   XOR2_X1 i_929 (.A(n_5310), .B(n_1025), .Z(n_1024));
   XOR2_X1 i_930 (.A(n_5290), .B(n_1026), .Z(n_1025));
   XNOR2_X1 i_931 (.A(n_1031), .B(n_1028), .ZN(n_1026));
   INV_X1 i_932 (.A(n_1028), .ZN(n_1027));
   AOI21_X1 i_933 (.A(n_1204), .B1(n_1279), .B2(n_1208), .ZN(n_1028));
   OAI21_X1 i_934 (.A(n_1032), .B1(n_1035), .B2(n_1033), .ZN(n_1031));
   NAND2_X1 i_935 (.A1(n_1035), .A2(n_1033), .ZN(n_1032));
   AND2_X1 i_936 (.A1(inputB[13]), .A2(inputA[30]), .ZN(n_1033));
   NAND2_X1 i_937 (.A1(inputB[12]), .A2(inputA[31]), .ZN(n_1035));
   INV_X1 i_938 (.A(n_1036), .ZN(n_5213));
   AOI21_X1 i_939 (.A(n_5210), .B1(n_5209), .B2(n_1116), .ZN(n_1036));
   INV_X1 i_940 (.A(n_1037), .ZN(n_5208));
   AOI21_X1 i_941 (.A(n_5205), .B1(n_5204), .B2(n_1119), .ZN(n_1037));
   XOR2_X1 i_942 (.A(n_5305), .B(n_1038), .Z(n_5307));
   XOR2_X1 i_943 (.A(n_5280), .B(n_1041), .Z(n_1038));
   NAND2_X1 i_944 (.A1(n_1193), .A2(n_1042), .ZN(n_1041));
   NAND2_X1 i_945 (.A1(n_1191), .A2(n_1189), .ZN(n_1042));
   INV_X1 i_946 (.A(n_1043), .ZN(n_5203));
   AOI21_X1 i_947 (.A(n_5200), .B1(n_5199), .B2(n_1134), .ZN(n_1043));
   XOR2_X1 i_948 (.A(n_5295), .B(n_1044), .Z(n_5297));
   XOR2_X1 i_949 (.A(n_1048), .B(n_1047), .Z(n_1044));
   NAND2_X1 i_950 (.A1(inputB[22]), .A2(inputA[21]), .ZN(n_1047));
   NAND2_X1 i_951 (.A1(n_1051), .A2(n_1049), .ZN(n_1048));
   INV_X1 i_952 (.A(n_1050), .ZN(n_1049));
   AOI22_X1 i_953 (.A1(inputB[21]), .A2(inputA[22]), .B1(inputB[20]), .B2(
      inputA[23]), .ZN(n_1050));
   NAND2_X1 i_954 (.A1(n_1194), .A2(n_1054), .ZN(n_1051));
   AND2_X1 i_955 (.A1(inputB[21]), .A2(inputA[23]), .ZN(n_1054));
   INV_X1 i_956 (.A(n_1055), .ZN(n_5193));
   AOI21_X1 i_957 (.A(n_5190), .B1(n_5189), .B2(n_1142), .ZN(n_1055));
   INV_X1 i_958 (.A(n_1057), .ZN(n_5198));
   AOI21_X1 i_959 (.A(n_5195), .B1(n_5194), .B2(n_1117), .ZN(n_1057));
   INV_X1 i_960 (.A(n_1058), .ZN(n_5183));
   AOI21_X1 i_961 (.A(n_5180), .B1(n_5179), .B2(n_1120), .ZN(n_1058));
   INV_X1 i_962 (.A(n_1059), .ZN(n_5188));
   AOI21_X1 i_963 (.A(n_5185), .B1(n_5184), .B2(n_1144), .ZN(n_1059));
   XOR2_X1 i_964 (.A(n_5285), .B(n_1060), .Z(n_5287));
   NAND2_X1 i_965 (.A1(n_1180), .A2(n_1061), .ZN(n_1060));
   NAND2_X1 i_966 (.A1(n_1177), .A2(n_1172), .ZN(n_1061));
   INV_X1 i_967 (.A(n_1062), .ZN(n_5178));
   AOI21_X1 i_968 (.A(n_5175), .B1(n_5174), .B2(n_1155), .ZN(n_1062));
   XOR2_X1 i_969 (.A(n_1064), .B(n_1063), .Z(n_5239));
   AND2_X1 i_970 (.A1(inputB[28]), .A2(inputA[15]), .ZN(n_1063));
   AND2_X1 i_971 (.A1(n_1066), .A2(n_1065), .ZN(n_1064));
   NAND2_X1 i_972 (.A1(n_1152), .A2(n_1071), .ZN(n_1065));
   NAND2_X1 i_973 (.A1(n_1151), .A2(n_1067), .ZN(n_1066));
   INV_X1 i_974 (.A(n_1071), .ZN(n_1067));
   NAND2_X1 i_975 (.A1(inputB[26]), .A2(inputA[17]), .ZN(n_1071));
   XOR2_X1 i_976 (.A(n_1076), .B(n_1075), .Z(n_5246));
   NAND2_X1 i_977 (.A1(inputB[25]), .A2(inputA[18]), .ZN(n_1075));
   NAND2_X1 i_978 (.A1(n_1082), .A2(n_1079), .ZN(n_1076));
   NAND2_X1 i_979 (.A1(n_1187), .A2(n_1080), .ZN(n_1079));
   INV_X1 i_980 (.A(n_1081), .ZN(n_1080));
   NAND2_X1 i_981 (.A1(inputB[24]), .A2(inputA[20]), .ZN(n_1081));
   INV_X1 i_982 (.A(n_1083), .ZN(n_1082));
   AOI22_X1 i_983 (.A1(inputB[24]), .A2(inputA[19]), .B1(inputB[23]), .B2(
      inputA[20]), .ZN(n_1083));
   XOR2_X1 i_984 (.A(n_1086), .B(n_1085), .Z(n_5260));
   AND2_X1 i_985 (.A1(inputB[19]), .A2(inputA[24]), .ZN(n_1085));
   AND2_X1 i_986 (.A1(n_1088), .A2(n_1087), .ZN(n_1086));
   NAND2_X1 i_987 (.A1(n_1129), .A2(n_1089), .ZN(n_1087));
   OR2_X1 i_988 (.A1(n_1129), .A2(n_1089), .ZN(n_1088));
   NAND2_X1 i_989 (.A1(inputB[17]), .A2(inputA[26]), .ZN(n_1089));
   XOR2_X1 i_990 (.A(n_1091), .B(n_1090), .Z(n_5267));
   NAND2_X1 i_991 (.A1(inputB[16]), .A2(inputA[27]), .ZN(n_1090));
   NAND2_X1 i_992 (.A1(n_1095), .A2(n_1093), .ZN(n_1091));
   INV_X1 i_993 (.A(n_1094), .ZN(n_1093));
   AOI22_X1 i_994 (.A1(inputB[15]), .A2(inputA[28]), .B1(inputB[14]), .B2(
      inputA[29]), .ZN(n_1094));
   NAND2_X1 i_995 (.A1(n_1201), .A2(n_1096), .ZN(n_1095));
   INV_X1 i_996 (.A(n_1100), .ZN(n_1096));
   NAND2_X1 i_997 (.A1(inputB[15]), .A2(inputA[29]), .ZN(n_1100));
   INV_X1 i_998 (.A(n_1104), .ZN(n_5168));
   AOI21_X1 i_999 (.A(n_5165), .B1(n_5164), .B2(n_1162), .ZN(n_1104));
   INV_X1 i_1000 (.A(n_1105), .ZN(n_5173));
   AOI21_X1 i_1001 (.A(n_5170), .B1(n_5169), .B2(n_1143), .ZN(n_1105));
   OAI21_X1 i_1002 (.A(n_1150), .B1(n_1149), .B2(n_1145), .ZN(n_5124));
   AOI22_X1 i_1003 (.A1(n_1298), .A2(n_1188), .B1(n_1185), .B2(n_1183), .ZN(
      n_5131));
   OAI21_X1 i_1004 (.A(n_1125), .B1(n_1124), .B2(n_1121), .ZN(n_5145));
   OAI21_X1 i_1005 (.A(n_1198), .B1(n_1200), .B2(n_1196), .ZN(n_5152));
   INV_X1 i_1006 (.A(n_1108), .ZN(n_5107));
   AOI21_X1 i_1007 (.A(n_5104), .B1(n_5103), .B2(n_1109), .ZN(n_1108));
   XNOR2_X1 i_1008 (.A(n_5093), .B(n_1115), .ZN(n_1109));
   XNOR2_X1 i_1009 (.A(n_5214), .B(n_1111), .ZN(n_5216));
   INV_X1 i_1010 (.A(n_1111), .ZN(n_1110));
   AOI21_X1 i_1011 (.A(n_5094), .B1(n_5093), .B2(n_1112), .ZN(n_1111));
   INV_X1 i_1012 (.A(n_1115), .ZN(n_1112));
   AOI21_X1 i_1013 (.A(n_4964), .B1(n_4963), .B2(n_1346), .ZN(n_1115));
   XOR2_X1 i_1014 (.A(n_5209), .B(n_1116), .Z(n_5211));
   XNOR2_X1 i_1015 (.A(n_5194), .B(n_1118), .ZN(n_1116));
   INV_X1 i_1016 (.A(n_1118), .ZN(n_1117));
   AOI21_X1 i_1017 (.A(n_5064), .B1(n_5063), .B2(n_1236), .ZN(n_1118));
   XOR2_X1 i_1018 (.A(n_5204), .B(n_1119), .Z(n_5206));
   XOR2_X1 i_1019 (.A(n_5179), .B(n_1120), .Z(n_1119));
   XOR2_X1 i_1020 (.A(n_1122), .B(n_1121), .Z(n_1120));
   NAND2_X1 i_1021 (.A1(inputB[19]), .A2(inputA[23]), .ZN(n_1121));
   NAND2_X1 i_1022 (.A1(n_1125), .A2(n_1123), .ZN(n_1122));
   INV_X1 i_1023 (.A(n_1124), .ZN(n_1123));
   AOI22_X1 i_1024 (.A1(inputB[18]), .A2(inputA[24]), .B1(inputB[17]), .B2(
      inputA[25]), .ZN(n_1124));
   NAND3_X1 i_1025 (.A1(inputB[18]), .A2(inputA[25]), .A3(n_1319), .ZN(n_1125));
   NAND2_X1 i_1026 (.A1(inputB[18]), .A2(inputA[25]), .ZN(n_1129));
   XNOR2_X1 i_1027 (.A(n_5199), .B(n_1138), .ZN(n_5201));
   INV_X1 i_1028 (.A(n_1138), .ZN(n_1134));
   AOI21_X1 i_1029 (.A(n_5079), .B1(n_5078), .B2(n_1234), .ZN(n_1138));
   INV_X1 i_1030 (.A(n_1139), .ZN(n_5092));
   AOI21_X1 i_1031 (.A(n_5089), .B1(n_5088), .B2(n_1226), .ZN(n_1139));
   INV_X1 i_1032 (.A(n_1140), .ZN(n_5087));
   AOI21_X1 i_1033 (.A(n_5084), .B1(n_5083), .B2(n_1228), .ZN(n_1140));
   XOR2_X1 i_1034 (.A(n_5189), .B(n_1142), .Z(n_5191));
   XOR2_X1 i_1035 (.A(n_5169), .B(n_1143), .Z(n_1142));
   AOI22_X1 i_1036 (.A1(n_1405), .A2(n_1292), .B1(n_1290), .B2(n_1288), .ZN(
      n_1143));
   XOR2_X1 i_1037 (.A(n_5184), .B(n_1144), .Z(n_5186));
   XOR2_X1 i_1038 (.A(n_1146), .B(n_1145), .Z(n_1144));
   NAND2_X1 i_1039 (.A1(inputB[28]), .A2(inputA[14]), .ZN(n_1145));
   NAND2_X1 i_1040 (.A1(n_1150), .A2(n_1148), .ZN(n_1146));
   INV_X1 i_1041 (.A(n_1149), .ZN(n_1148));
   AOI22_X1 i_1042 (.A1(inputB[27]), .A2(inputA[15]), .B1(inputB[26]), .B2(
      inputA[16]), .ZN(n_1149));
   NAND2_X1 i_1043 (.A1(n_1291), .A2(n_1151), .ZN(n_1150));
   INV_X1 i_1044 (.A(n_1152), .ZN(n_1151));
   NAND2_X1 i_1045 (.A1(inputB[27]), .A2(inputA[16]), .ZN(n_1152));
   INV_X1 i_1046 (.A(n_1153), .ZN(n_5077));
   AOI21_X1 i_1047 (.A(n_5074), .B1(n_5073), .B2(n_1231), .ZN(n_1153));
   XNOR2_X1 i_1048 (.A(n_5174), .B(n_1156), .ZN(n_5176));
   INV_X1 i_1049 (.A(n_1156), .ZN(n_1155));
   AOI21_X1 i_1050 (.A(n_5044), .B1(n_5043), .B2(n_1284), .ZN(n_1156));
   INV_X1 i_1051 (.A(n_1157), .ZN(n_5062));
   AOI21_X1 i_1053 (.A(n_5059), .B1(n_5058), .B2(n_1265), .ZN(n_1157));
   INV_X1 i_1054 (.A(n_1158), .ZN(n_5072));
   AOI21_X1 i_1055 (.A(n_5069), .B1(n_5068), .B2(n_1248), .ZN(n_1158));
   XOR2_X1 i_1056 (.A(n_5164), .B(n_1162), .Z(n_5166));
   OAI21_X1 i_1057 (.A(n_1309), .B1(n_1318), .B2(n_1304), .ZN(n_1162));
   INV_X1 i_1058 (.A(n_1167), .ZN(n_5057));
   AOI21_X1 i_1059 (.A(n_5054), .B1(n_5053), .B2(n_1285), .ZN(n_1167));
   XOR2_X1 i_1060 (.A(n_1176), .B(n_1172), .Z(n_5114));
   NAND2_X1 i_1061 (.A1(inputB[31]), .A2(inputA[11]), .ZN(n_1172));
   AND2_X1 i_1062 (.A1(n_1180), .A2(n_1177), .ZN(n_1176));
   NAND2_X1 i_1063 (.A1(n_1259), .A2(n_1182), .ZN(n_1177));
   NAND2_X1 i_1064 (.A1(n_1255), .A2(n_1181), .ZN(n_1180));
   INV_X1 i_1065 (.A(n_1182), .ZN(n_1181));
   NAND2_X1 i_1066 (.A1(inputB[29]), .A2(inputA[13]), .ZN(n_1182));
   XOR2_X1 i_1068 (.A(n_1184), .B(n_1183), .Z(n_5130));
   NAND2_X1 i_1069 (.A1(inputB[25]), .A2(inputA[17]), .ZN(n_1183));
   OAI21_X1 i_1070 (.A(n_1185), .B1(n_1297), .B2(n_1187), .ZN(n_1184));
   NAND2_X1 i_1072 (.A1(n_1297), .A2(n_1187), .ZN(n_1185));
   INV_X1 i_1073 (.A(n_1188), .ZN(n_1187));
   NAND2_X1 i_1074 (.A1(inputB[23]), .A2(inputA[19]), .ZN(n_1188));
   XOR2_X1 i_1075 (.A(n_1190), .B(n_1189), .Z(n_5137));
   AND2_X1 i_1076 (.A1(inputB[22]), .A2(inputA[20]), .ZN(n_1189));
   AND2_X1 i_1077 (.A1(n_1193), .A2(n_1191), .ZN(n_1190));
   NAND2_X1 i_1078 (.A1(n_1247), .A2(n_1195), .ZN(n_1191));
   NAND2_X1 i_1079 (.A1(n_1246), .A2(n_1194), .ZN(n_1193));
   INV_X1 i_1080 (.A(n_1195), .ZN(n_1194));
   NAND2_X1 i_1081 (.A1(inputB[20]), .A2(inputA[22]), .ZN(n_1195));
   XOR2_X1 i_1082 (.A(n_1197), .B(n_1196), .Z(n_5151));
   NAND2_X1 i_1083 (.A1(inputB[16]), .A2(inputA[26]), .ZN(n_1196));
   NAND2_X1 i_1084 (.A1(n_1199), .A2(n_1198), .ZN(n_1197));
   NAND3_X1 i_1085 (.A1(inputB[15]), .A2(inputA[27]), .A3(n_1201), .ZN(n_1198));
   INV_X1 i_1086 (.A(n_1200), .ZN(n_1199));
   AOI21_X1 i_1087 (.A(n_1201), .B1(inputB[15]), .B2(inputA[27]), .ZN(n_1200));
   AND2_X1 i_1088 (.A1(inputB[14]), .A2(inputA[28]), .ZN(n_1201));
   XOR2_X1 i_1089 (.A(n_1279), .B(n_1202), .Z(n_5157));
   NAND2_X1 i_1090 (.A1(n_1208), .A2(n_1203), .ZN(n_1202));
   INV_X1 i_1091 (.A(n_1204), .ZN(n_1203));
   AOI211_X1 i_1092 (.A(n_5758), .B(n_5753), .C1(inputB[13]), .C2(inputA[29]), 
      .ZN(n_1204));
   OAI211_X1 i_1093 (.A(inputB[13]), .B(inputA[29]), .C1(n_5758), .C2(n_5753), 
      .ZN(n_1208));
   INV_X1 i_1095 (.A(n_1209), .ZN(n_5052));
   AOI21_X1 i_1096 (.A(n_5049), .B1(n_5048), .B2(n_1233), .ZN(n_1209));
   AOI21_X1 i_1097 (.A(n_1263), .B1(n_1264), .B2(n_1254), .ZN(n_4995));
   OAI21_X1 i_1099 (.A(n_1295), .B1(n_1300), .B2(n_1293), .ZN(n_5011));
   OAI21_X1 i_1100 (.A(n_1243), .B1(n_1242), .B2(n_1237), .ZN(n_5018));
   OAI21_X1 i_1101 (.A(n_1329), .B1(n_1332), .B2(n_1324), .ZN(n_5032));
   OAI21_X1 i_1102 (.A(n_1278), .B1(n_1277), .B2(n_1269), .ZN(n_5039));
   INV_X1 i_1103 (.A(n_1212), .ZN(n_4987));
   AOI21_X1 i_1104 (.A(n_4984), .B1(n_4983), .B2(n_1213), .ZN(n_1212));
   INV_X1 i_1105 (.A(n_1218), .ZN(n_1213));
   AOI21_X1 i_1106 (.A(n_4851), .B1(n_4850), .B2(n_1465), .ZN(n_1218));
   XNOR2_X1 i_1107 (.A(n_5098), .B(n_1223), .ZN(n_5100));
   INV_X1 i_1108 (.A(n_1223), .ZN(n_1222));
   AOI21_X1 i_1109 (.A(n_4974), .B1(n_4973), .B2(n_1340), .ZN(n_1223));
   INV_X1 i_1110 (.A(n_1225), .ZN(n_4982));
   AOI21_X1 i_1111 (.A(n_4979), .B1(n_4978), .B2(n_1337), .ZN(n_1225));
   XNOR2_X1 i_1112 (.A(n_5088), .B(n_1227), .ZN(n_5090));
   INV_X1 i_1113 (.A(n_1227), .ZN(n_1226));
   AOI21_X1 i_1114 (.A(n_4959), .B1(n_4958), .B2(n_1353), .ZN(n_1227));
   XNOR2_X1 i_1115 (.A(n_5083), .B(n_1229), .ZN(n_5085));
   INV_X1 i_1116 (.A(n_1229), .ZN(n_1228));
   AOI21_X1 i_1117 (.A(n_4954), .B1(n_4953), .B2(n_1350), .ZN(n_1229));
   INV_X1 i_1118 (.A(n_1230), .ZN(n_4972));
   AOI21_X1 i_1119 (.A(n_4969), .B1(n_4968), .B2(n_1342), .ZN(n_1230));
   XOR2_X1 i_1120 (.A(n_5073), .B(n_1231), .Z(n_5075));
   XOR2_X1 i_1122 (.A(n_5048), .B(n_1233), .Z(n_1231));
   AOI21_X1 i_1123 (.A(n_1377), .B1(n_1381), .B2(n_1371), .ZN(n_1233));
   XNOR2_X1 i_1124 (.A(n_5078), .B(n_1235), .ZN(n_5080));
   INV_X1 i_1126 (.A(n_1235), .ZN(n_1234));
   AOI21_X1 i_1127 (.A(n_4939), .B1(n_4938), .B2(n_1356), .ZN(n_1235));
   XOR2_X1 i_1128 (.A(n_5063), .B(n_1236), .Z(n_5065));
   XOR2_X1 i_1130 (.A(n_1240), .B(n_1237), .Z(n_1236));
   NAND2_X1 i_1131 (.A1(inputB[22]), .A2(inputA[19]), .ZN(n_1237));
   NAND2_X1 i_1132 (.A1(n_1243), .A2(n_1241), .ZN(n_1240));
   INV_X1 i_1133 (.A(n_1242), .ZN(n_1241));
   AOI22_X1 i_1134 (.A1(inputB[21]), .A2(inputA[20]), .B1(inputB[20]), .B2(
      inputA[21]), .ZN(n_1242));
   NAND2_X1 i_1135 (.A1(n_1413), .A2(n_1246), .ZN(n_1243));
   INV_X1 i_1136 (.A(n_1247), .ZN(n_1246));
   NAND2_X1 i_1137 (.A1(inputB[21]), .A2(inputA[21]), .ZN(n_1247));
   XOR2_X1 i_1138 (.A(n_5068), .B(n_1248), .Z(n_5070));
   XNOR2_X1 i_1139 (.A(n_1264), .B(n_1249), .ZN(n_1248));
   NOR2_X1 i_1140 (.A1(n_1263), .A2(n_1250), .ZN(n_1249));
   INV_X1 i_1141 (.A(n_1254), .ZN(n_1250));
   NAND3_X1 i_1142 (.A1(inputB[29]), .A2(inputA[11]), .A3(n_1255), .ZN(n_1254));
   INV_X1 i_1143 (.A(n_1259), .ZN(n_1255));
   NAND2_X1 i_1144 (.A1(inputB[30]), .A2(inputA[12]), .ZN(n_1259));
   AOI22_X1 i_1145 (.A1(inputB[30]), .A2(inputA[11]), .B1(inputB[29]), .B2(
      inputA[12]), .ZN(n_1263));
   AND2_X1 i_1146 (.A1(inputB[31]), .A2(inputA[10]), .ZN(n_1264));
   XOR2_X1 i_1147 (.A(n_5058), .B(n_1265), .Z(n_5060));
   XOR2_X1 i_1148 (.A(n_1273), .B(n_1269), .Z(n_1265));
   NAND2_X1 i_1149 (.A1(inputB[13]), .A2(inputA[28]), .ZN(n_1269));
   NAND2_X1 i_1150 (.A1(n_1278), .A2(n_1274), .ZN(n_1273));
   INV_X1 i_1152 (.A(n_1277), .ZN(n_1274));
   AOI22_X1 i_1153 (.A1(inputB[12]), .A2(inputA[29]), .B1(inputB[11]), .B2(
      inputA[30]), .ZN(n_1277));
   NAND3_X1 i_1154 (.A1(inputB[12]), .A2(inputA[30]), .A3(n_1430), .ZN(n_1278));
   NAND2_X1 i_1156 (.A1(inputB[12]), .A2(inputA[30]), .ZN(n_1279));
   INV_X1 i_1157 (.A(n_1280), .ZN(n_4952));
   AOI21_X1 i_1158 (.A(n_4949), .B1(n_4948), .B2(n_1347), .ZN(n_1280));
   INV_X1 i_1160 (.A(n_1281), .ZN(n_4947));
   AOI21_X1 i_1161 (.A(n_4944), .B1(n_4943), .B2(n_1367), .ZN(n_1281));
   XOR2_X1 i_1162 (.A(n_5043), .B(n_1284), .Z(n_5045));
   OAI21_X1 i_1164 (.A(n_1360), .B1(n_1363), .B2(n_1357), .ZN(n_1284));
   XNOR2_X1 i_1165 (.A(n_5053), .B(n_1286), .ZN(n_5055));
   INV_X1 i_1166 (.A(n_1286), .ZN(n_1285));
   AOI21_X1 i_1167 (.A(n_4929), .B1(n_4928), .B2(n_1393), .ZN(n_1286));
   INV_X1 i_1168 (.A(n_1287), .ZN(n_4937));
   AOI21_X1 i_1169 (.A(n_4934), .B1(n_4933), .B2(n_1354), .ZN(n_1287));
   XOR2_X1 i_1170 (.A(n_1289), .B(n_1288), .Z(n_5003));
   NAND2_X1 i_1171 (.A1(inputB[28]), .A2(inputA[13]), .ZN(n_1288));
   OAI21_X1 i_1172 (.A(n_1290), .B1(n_1404), .B2(n_1291), .ZN(n_1289));
   NAND2_X1 i_1173 (.A1(n_1404), .A2(n_1291), .ZN(n_1290));
   INV_X1 i_1174 (.A(n_1292), .ZN(n_1291));
   NAND2_X1 i_1175 (.A1(inputB[26]), .A2(inputA[15]), .ZN(n_1292));
   XOR2_X1 i_1176 (.A(n_1294), .B(n_1293), .Z(n_5010));
   NAND2_X1 i_1177 (.A1(inputB[25]), .A2(inputA[16]), .ZN(n_1293));
   NAND2_X1 i_1178 (.A1(n_1299), .A2(n_1295), .ZN(n_1294));
   NAND3_X1 i_1179 (.A1(inputB[23]), .A2(inputA[17]), .A3(n_1297), .ZN(n_1295));
   INV_X1 i_1180 (.A(n_1298), .ZN(n_1297));
   NAND2_X1 i_1181 (.A1(inputB[24]), .A2(inputA[18]), .ZN(n_1298));
   INV_X1 i_1182 (.A(n_1300), .ZN(n_1299));
   AOI22_X1 i_1183 (.A1(inputB[24]), .A2(inputA[17]), .B1(inputB[23]), .B2(
      inputA[18]), .ZN(n_1300));
   XOR2_X1 i_1184 (.A(n_1305), .B(n_1304), .Z(n_5024));
   NAND2_X1 i_1185 (.A1(inputB[19]), .A2(inputA[22]), .ZN(n_1304));
   NAND2_X1 i_1186 (.A1(n_1314), .A2(n_1309), .ZN(n_1305));
   NAND3_X1 i_1187 (.A1(inputB[18]), .A2(inputA[23]), .A3(n_1319), .ZN(n_1309));
   INV_X1 i_1188 (.A(n_1318), .ZN(n_1314));
   AOI21_X1 i_1189 (.A(n_1319), .B1(inputB[18]), .B2(inputA[23]), .ZN(n_1318));
   AND2_X1 i_1190 (.A1(inputB[17]), .A2(inputA[24]), .ZN(n_1319));
   XOR2_X1 i_1191 (.A(n_1328), .B(n_1324), .Z(n_5031));
   NAND2_X1 i_1192 (.A1(inputB[16]), .A2(inputA[25]), .ZN(n_1324));
   NAND2_X1 i_1194 (.A1(n_1331), .A2(n_1329), .ZN(n_1328));
   NAND3_X1 i_1195 (.A1(inputB[14]), .A2(inputA[27]), .A3(n_1361), .ZN(n_1329));
   INV_X1 i_1196 (.A(n_1332), .ZN(n_1331));
   AOI21_X1 i_1198 (.A(n_1361), .B1(inputB[14]), .B2(inputA[27]), .ZN(n_1332));
   AOI21_X1 i_1199 (.A(n_1455), .B1(n_1450), .B2(n_1434), .ZN(n_4918));
   INV_X1 i_1200 (.A(n_1333), .ZN(n_4927));
   AOI21_X1 i_1202 (.A(n_4924), .B1(n_4923), .B2(n_1392), .ZN(n_1333));
   OAI21_X1 i_1203 (.A(n_1397), .B1(n_1399), .B2(n_1395), .ZN(n_4867));
   OAI21_X1 i_1204 (.A(n_1403), .B1(n_1409), .B2(n_1401), .ZN(n_4876));
   AOI22_X1 i_1206 (.A1(n_1557), .A2(n_1414), .B1(n_1412), .B2(n_1410), .ZN(
      n_4890));
   OAI21_X1 i_1207 (.A(n_1418), .B1(n_1421), .B2(n_1416), .ZN(n_4897));
   OAI21_X1 i_1208 (.A(n_1424), .B1(n_1426), .B2(n_1422), .ZN(n_4911));
   NAND2_X1 i_1209 (.A1(inputB[10]), .A2(inputA[31]), .ZN(n_382));
   INV_X1 i_1210 (.A(n_1334), .ZN(n_4859));
   AOI21_X1 i_1211 (.A(n_4856), .B1(n_4855), .B2(n_1335), .ZN(n_1334));
   INV_X1 i_1212 (.A(n_1336), .ZN(n_1335));
   AOI21_X1 i_1213 (.A(n_4718), .B1(n_4717), .B2(n_1577), .ZN(n_1336));
   XNOR2_X1 i_1214 (.A(n_4978), .B(n_1339), .ZN(n_4980));
   INV_X1 i_1215 (.A(n_1339), .ZN(n_1337));
   AOI21_X1 i_1216 (.A(n_4846), .B1(n_4845), .B2(n_1470), .ZN(n_1339));
   XNOR2_X1 i_1217 (.A(n_4973), .B(n_1341), .ZN(n_4975));
   INV_X1 i_1218 (.A(n_1341), .ZN(n_1340));
   AOI21_X1 i_1219 (.A(n_4836), .B1(n_4835), .B2(n_1481), .ZN(n_1341));
   XNOR2_X1 i_1220 (.A(n_4968), .B(n_1343), .ZN(n_4970));
   INV_X1 i_1221 (.A(n_1343), .ZN(n_1342));
   AOI21_X1 i_1222 (.A(n_4831), .B1(n_4830), .B2(n_1471), .ZN(n_1343));
   XOR2_X1 i_1223 (.A(n_4963), .B(n_1346), .Z(n_4965));
   XNOR2_X1 i_1224 (.A(n_4948), .B(n_1348), .ZN(n_1346));
   INV_X1 i_1225 (.A(n_1348), .ZN(n_1347));
   AOI21_X1 i_1226 (.A(n_4801), .B1(n_4800), .B2(n_1496), .ZN(n_1348));
   INV_X1 i_1227 (.A(n_1349), .ZN(n_4844));
   AOI21_X1 i_1228 (.A(n_4841), .B1(n_4840), .B2(n_1466), .ZN(n_1349));
   XNOR2_X1 i_1229 (.A(n_4953), .B(n_1352), .ZN(n_4955));
   INV_X1 i_1230 (.A(n_1352), .ZN(n_1350));
   AOI21_X1 i_1231 (.A(n_4816), .B1(n_4815), .B2(n_1483), .ZN(n_1352));
   XOR2_X1 i_1232 (.A(n_4958), .B(n_1353), .Z(n_4960));
   XNOR2_X1 i_1233 (.A(n_4933), .B(n_1355), .ZN(n_1353));
   INV_X1 i_1234 (.A(n_1355), .ZN(n_1354));
   AOI21_X1 i_1236 (.A(n_4791), .B1(n_4790), .B2(n_1533), .ZN(n_1355));
   XOR2_X1 i_1237 (.A(n_4938), .B(n_1356), .Z(n_4940));
   XOR2_X1 i_1238 (.A(n_1358), .B(n_1357), .Z(n_1356));
   NAND2_X1 i_1240 (.A1(inputB[16]), .A2(inputA[24]), .ZN(n_1357));
   NAND2_X1 i_1241 (.A1(n_1362), .A2(n_1360), .ZN(n_1358));
   NAND2_X1 i_1242 (.A1(n_1564), .A2(n_1361), .ZN(n_1360));
   AND2_X1 i_1244 (.A1(inputB[15]), .A2(inputA[26]), .ZN(n_1361));
   INV_X1 i_1245 (.A(n_1363), .ZN(n_1362));
   AOI22_X1 i_1246 (.A1(inputB[15]), .A2(inputA[25]), .B1(inputB[14]), .B2(
      inputA[26]), .ZN(n_1363));
   XOR2_X1 i_1248 (.A(n_4943), .B(n_1367), .Z(n_4945));
   XOR2_X1 i_1249 (.A(n_1372), .B(n_1371), .Z(n_1367));
   NAND2_X1 i_1250 (.A1(inputB[25]), .A2(inputA[15]), .ZN(n_1371));
   NAND2_X1 i_1252 (.A1(n_1381), .A2(n_1373), .ZN(n_1372));
   INV_X1 i_1253 (.A(n_1377), .ZN(n_1373));
   AOI22_X1 i_1254 (.A1(inputB[24]), .A2(inputA[16]), .B1(inputB[23]), .B2(
      inputA[17]), .ZN(n_1377));
   NAND3_X1 i_1255 (.A1(inputB[24]), .A2(inputA[17]), .A3(n_1551), .ZN(n_1381));
   INV_X1 i_1256 (.A(n_1382), .ZN(n_4824));
   AOI21_X1 i_1257 (.A(n_4821), .B1(n_4820), .B2(n_1493), .ZN(n_1382));
   INV_X1 i_1258 (.A(n_1387), .ZN(n_4829));
   AOI21_X1 i_1259 (.A(n_4826), .B1(n_4825), .B2(n_1491), .ZN(n_1387));
   INV_X1 i_1260 (.A(n_1388), .ZN(n_4809));
   AOI21_X1 i_1261 (.A(n_4806), .B1(n_4805), .B2(n_1472), .ZN(n_1388));
   INV_X1 i_1262 (.A(n_1391), .ZN(n_4814));
   AOI21_X1 i_1263 (.A(n_4811), .B1(n_4810), .B2(n_1501), .ZN(n_1391));
   XOR2_X1 i_1264 (.A(n_4923), .B(n_1392), .Z(n_4925));
   AOI21_X1 i_1265 (.A(n_1512), .B1(n_1517), .B2(n_1502), .ZN(n_1392));
   XOR2_X1 i_1266 (.A(n_4928), .B(n_1393), .Z(n_4930));
   OAI21_X1 i_1267 (.A(n_1486), .B1(n_1488), .B2(n_1484), .ZN(n_1393));
   XOR2_X1 i_1268 (.A(n_1396), .B(n_1395), .Z(n_4866));
   AND2_X1 i_1269 (.A1(inputB[31]), .A2(inputA[9]), .ZN(n_1395));
   NAND2_X1 i_1270 (.A1(n_1398), .A2(n_1397), .ZN(n_1396));
   NAND3_X1 i_1271 (.A1(inputB[30]), .A2(inputA[11]), .A3(n_1542), .ZN(n_1397));
   INV_X1 i_1272 (.A(n_1399), .ZN(n_1398));
   AOI22_X1 i_1273 (.A1(inputB[30]), .A2(inputA[10]), .B1(inputB[29]), .B2(
      inputA[11]), .ZN(n_1399));
   XOR2_X1 i_1274 (.A(n_1402), .B(n_1401), .Z(n_4875));
   NAND2_X1 i_1275 (.A1(inputB[28]), .A2(inputA[12]), .ZN(n_1401));
   NAND2_X1 i_1276 (.A1(n_1406), .A2(n_1403), .ZN(n_1402));
   NAND3_X1 i_1277 (.A1(inputB[26]), .A2(inputA[13]), .A3(n_1404), .ZN(n_1403));
   INV_X1 i_1278 (.A(n_1405), .ZN(n_1404));
   NAND2_X1 i_1279 (.A1(inputB[27]), .A2(inputA[14]), .ZN(n_1405));
   INV_X1 i_1281 (.A(n_1409), .ZN(n_1406));
   AOI22_X1 i_1282 (.A1(inputB[27]), .A2(inputA[13]), .B1(inputB[26]), .B2(
      inputA[14]), .ZN(n_1409));
   XOR2_X1 i_1283 (.A(n_1411), .B(n_1410), .Z(n_4889));
   NAND2_X1 i_1285 (.A1(inputB[22]), .A2(inputA[18]), .ZN(n_1410));
   OAI21_X1 i_1286 (.A(n_1412), .B1(n_1556), .B2(n_1413), .ZN(n_1411));
   NAND2_X1 i_1287 (.A1(n_1556), .A2(n_1413), .ZN(n_1412));
   INV_X1 i_1289 (.A(n_1414), .ZN(n_1413));
   NAND2_X1 i_1290 (.A1(inputB[20]), .A2(inputA[20]), .ZN(n_1414));
   XOR2_X1 i_1291 (.A(n_1417), .B(n_1416), .Z(n_4896));
   NAND2_X1 i_1293 (.A1(inputB[19]), .A2(inputA[21]), .ZN(n_1416));
   NAND2_X1 i_1294 (.A1(n_1419), .A2(n_1418), .ZN(n_1417));
   NAND3_X1 i_1295 (.A1(inputB[17]), .A2(inputA[23]), .A3(n_1521), .ZN(n_1418));
   INV_X1 i_1297 (.A(n_1421), .ZN(n_1419));
   AOI21_X1 i_1298 (.A(n_1521), .B1(inputB[17]), .B2(inputA[23]), .ZN(n_1421));
   XOR2_X1 i_1299 (.A(n_1423), .B(n_1422), .Z(n_4910));
   NAND2_X1 i_1301 (.A1(inputB[13]), .A2(inputA[27]), .ZN(n_1422));
   NAND2_X1 i_1302 (.A1(n_1425), .A2(n_1424), .ZN(n_1423));
   NAND3_X1 i_1303 (.A1(inputB[12]), .A2(inputA[28]), .A3(n_1430), .ZN(n_1424));
   INV_X1 i_1304 (.A(n_1426), .ZN(n_1425));
   AOI21_X1 i_1305 (.A(n_1430), .B1(inputB[12]), .B2(inputA[28]), .ZN(n_1426));
   NOR2_X1 i_1306 (.A1(n_5758), .A2(n_5750), .ZN(n_1430));
   XOR2_X1 i_1307 (.A(n_1440), .B(n_1435), .Z(n_4917));
   INV_X1 i_1308 (.A(n_1435), .ZN(n_1434));
   AOI21_X1 i_1309 (.A(n_1478), .B1(n_1475), .B2(n_1473), .ZN(n_1435));
   NOR2_X1 i_1310 (.A1(n_1455), .A2(n_1445), .ZN(n_1440));
   INV_X1 i_1311 (.A(n_1450), .ZN(n_1445));
   OAI211_X1 i_1312 (.A(inputB[10]), .B(inputA[30]), .C1(n_5757), .C2(n_5753), 
      .ZN(n_1450));
   AOI211_X1 i_1313 (.A(n_5757), .B(n_5753), .C1(inputB[10]), .C2(inputA[30]), 
      .ZN(n_1455));
   INV_X1 i_1314 (.A(n_1459), .ZN(n_4799));
   AOI21_X1 i_1315 (.A(n_4796), .B1(n_4795), .B2(n_1535), .ZN(n_1459));
   NAND2_X1 i_1316 (.A1(n_1541), .A2(n_1460), .ZN(n_4734));
   NAND2_X1 i_1317 (.A1(n_1539), .A2(n_1537), .ZN(n_1460));
   OAI21_X1 i_1318 (.A(n_1546), .B1(n_1550), .B2(n_1544), .ZN(n_4750));
   OAI21_X1 i_1319 (.A(n_1554), .B1(n_1559), .B2(n_1552), .ZN(n_4757));
   AOI22_X1 i_1320 (.A1(n_1631), .A2(n_1565), .B1(n_1563), .B2(n_1560), .ZN(
      n_4771));
   OAI21_X1 i_1321 (.A(n_1568), .B1(n_1570), .B2(n_1566), .ZN(n_4778));
   INV_X1 i_1322 (.A(n_1462), .ZN(n_4726));
   AOI21_X1 i_1323 (.A(n_4723), .B1(n_4722), .B2(n_1463), .ZN(n_1462));
   INV_X1 i_1324 (.A(n_1464), .ZN(n_1463));
   AOI21_X1 i_1325 (.A(n_4581), .B1(n_4580), .B2(n_1721), .ZN(n_1464));
   XOR2_X1 i_1326 (.A(n_4850), .B(n_1465), .Z(n_4852));
   XNOR2_X1 i_1327 (.A(n_4840), .B(n_1467), .ZN(n_1465));
   INV_X1 i_1328 (.A(n_1467), .ZN(n_1466));
   AOI21_X1 i_1329 (.A(n_4698), .B1(n_4697), .B2(n_1598), .ZN(n_1467));
   XOR2_X1 i_1330 (.A(n_4845), .B(n_1470), .Z(n_4847));
   XOR2_X1 i_1331 (.A(n_4830), .B(n_1471), .Z(n_1470));
   XOR2_X1 i_1332 (.A(n_4805), .B(n_1472), .Z(n_1471));
   XNOR2_X1 i_1333 (.A(n_1474), .B(n_1473), .ZN(n_1472));
   NAND2_X1 i_1334 (.A1(inputB[10]), .A2(inputA[29]), .ZN(n_1473));
   NOR2_X1 i_1335 (.A1(n_1478), .A2(n_1477), .ZN(n_1474));
   INV_X1 i_1336 (.A(n_1477), .ZN(n_1475));
   AOI21_X1 i_1338 (.A(n_1714), .B1(inputB[8]), .B2(inputA[31]), .ZN(n_1477));
   AND3_X1 i_1339 (.A1(inputB[8]), .A2(inputA[31]), .A3(n_1714), .ZN(n_1478));
   INV_X1 i_1340 (.A(n_1479), .ZN(n_4716));
   AOI21_X1 i_1342 (.A(n_4713), .B1(n_4712), .B2(n_1597), .ZN(n_1479));
   INV_X1 i_1343 (.A(n_1480), .ZN(n_4711));
   AOI21_X1 i_1344 (.A(n_4708), .B1(n_4707), .B2(n_1582), .ZN(n_1480));
   XOR2_X1 i_1346 (.A(n_4835), .B(n_1481), .Z(n_4837));
   XOR2_X1 i_1347 (.A(n_4815), .B(n_1483), .Z(n_1481));
   XOR2_X1 i_1348 (.A(n_1485), .B(n_1484), .Z(n_1483));
   NAND2_X1 i_1350 (.A1(inputB[28]), .A2(inputA[11]), .ZN(n_1484));
   NAND2_X1 i_1351 (.A1(n_1487), .A2(n_1486), .ZN(n_1485));
   NAND4_X1 i_1352 (.A1(inputB[26]), .A2(inputA[12]), .A3(inputB[27]), .A4(
      inputA[13]), .ZN(n_1486));
   INV_X1 i_1354 (.A(n_1488), .ZN(n_1487));
   AOI22_X1 i_1355 (.A1(inputB[27]), .A2(inputA[12]), .B1(inputB[26]), .B2(
      inputA[13]), .ZN(n_1488));
   INV_X1 i_1356 (.A(n_1490), .ZN(n_4706));
   AOI21_X1 i_1358 (.A(n_4703), .B1(n_4702), .B2(n_1607), .ZN(n_1490));
   XNOR2_X1 i_1359 (.A(n_4825), .B(n_1492), .ZN(n_4827));
   INV_X1 i_1360 (.A(n_1492), .ZN(n_1491));
   AOI21_X1 i_1361 (.A(n_4678), .B1(n_4677), .B2(n_1611), .ZN(n_1492));
   XOR2_X1 i_1362 (.A(n_4820), .B(n_1493), .Z(n_4822));
   XNOR2_X1 i_1363 (.A(n_4800), .B(n_1497), .ZN(n_1493));
   INV_X1 i_1364 (.A(n_1497), .ZN(n_1496));
   AOI21_X1 i_1365 (.A(n_4663), .B1(n_4662), .B2(n_1649), .ZN(n_1497));
   XOR2_X1 i_1366 (.A(n_4810), .B(n_1501), .Z(n_4812));
   XOR2_X1 i_1367 (.A(n_1506), .B(n_1502), .Z(n_1501));
   NAND2_X1 i_1368 (.A1(inputB[19]), .A2(inputA[20]), .ZN(n_1502));
   NAND2_X1 i_1369 (.A1(n_1517), .A2(n_1507), .ZN(n_1506));
   INV_X1 i_1370 (.A(n_1512), .ZN(n_1507));
   AOI22_X1 i_1371 (.A1(inputB[18]), .A2(inputA[21]), .B1(inputB[17]), .B2(
      inputA[22]), .ZN(n_1512));
   NAND2_X1 i_1372 (.A1(n_1703), .A2(n_1521), .ZN(n_1517));
   AND2_X1 i_1373 (.A1(inputB[18]), .A2(inputA[22]), .ZN(n_1521));
   INV_X1 i_1374 (.A(n_1522), .ZN(n_4691));
   AOI21_X1 i_1375 (.A(n_4688), .B1(n_4687), .B2(n_1622), .ZN(n_1522));
   INV_X1 i_1376 (.A(n_1527), .ZN(n_4696));
   AOI21_X1 i_1377 (.A(n_4693), .B1(n_4692), .B2(n_1583), .ZN(n_1527));
   INV_X1 i_1378 (.A(n_1531), .ZN(n_4686));
   AOI21_X1 i_1379 (.A(n_4683), .B1(n_4682), .B2(n_1634), .ZN(n_1531));
   INV_X1 i_1380 (.A(n_1532), .ZN(n_4676));
   AOI21_X1 i_1381 (.A(n_4673), .B1(n_4672), .B2(n_1625), .ZN(n_1532));
   XOR2_X1 i_1382 (.A(n_4790), .B(n_1533), .Z(n_4792));
   OAI21_X1 i_1383 (.A(n_1629), .B1(n_1633), .B2(n_1626), .ZN(n_1533));
   XOR2_X1 i_1384 (.A(n_4795), .B(n_1535), .Z(n_4797));
   OAI21_X1 i_1385 (.A(n_1615), .B1(n_1617), .B2(n_1612), .ZN(n_1535));
   INV_X1 i_1386 (.A(n_1536), .ZN(n_4671));
   AOI21_X1 i_1387 (.A(n_4668), .B1(n_4667), .B2(n_1638), .ZN(n_1536));
   XOR2_X1 i_1388 (.A(n_1538), .B(n_1537), .Z(n_4733));
   NAND2_X1 i_1389 (.A1(inputB[31]), .A2(inputA[8]), .ZN(n_1537));
   AND2_X1 i_1390 (.A1(n_1541), .A2(n_1539), .ZN(n_1538));
   NAND2_X1 i_1391 (.A1(n_1658), .A2(n_1543), .ZN(n_1539));
   NAND2_X1 i_1392 (.A1(n_1657), .A2(n_1542), .ZN(n_1541));
   INV_X1 i_1393 (.A(n_1543), .ZN(n_1542));
   NAND2_X1 i_1395 (.A1(inputB[29]), .A2(inputA[10]), .ZN(n_1543));
   XOR2_X1 i_1396 (.A(n_1545), .B(n_1544), .Z(n_4749));
   NAND2_X1 i_1397 (.A1(inputB[25]), .A2(inputA[14]), .ZN(n_1544));
   NAND2_X1 i_1399 (.A1(n_1549), .A2(n_1546), .ZN(n_1545));
   NAND3_X1 i_1400 (.A1(inputB[24]), .A2(inputA[15]), .A3(n_1551), .ZN(n_1546));
   INV_X1 i_1401 (.A(n_1550), .ZN(n_1549));
   AOI21_X1 i_1403 (.A(n_1551), .B1(inputB[24]), .B2(inputA[15]), .ZN(n_1550));
   AND2_X1 i_1404 (.A1(inputB[23]), .A2(inputA[16]), .ZN(n_1551));
   XOR2_X1 i_1405 (.A(n_1553), .B(n_1552), .Z(n_4756));
   NAND2_X1 i_1407 (.A1(inputB[22]), .A2(inputA[17]), .ZN(n_1552));
   NAND2_X1 i_1408 (.A1(n_1558), .A2(n_1554), .ZN(n_1553));
   NAND2_X1 i_1409 (.A1(n_1692), .A2(n_1556), .ZN(n_1554));
   INV_X1 i_1411 (.A(n_1557), .ZN(n_1556));
   NAND2_X1 i_1412 (.A1(inputB[21]), .A2(inputA[19]), .ZN(n_1557));
   INV_X1 i_1413 (.A(n_1559), .ZN(n_1558));
   AOI22_X1 i_1415 (.A1(inputB[21]), .A2(inputA[18]), .B1(inputB[20]), .B2(
      inputA[19]), .ZN(n_1559));
   XOR2_X1 i_1416 (.A(n_1562), .B(n_1560), .Z(n_4770));
   NAND2_X1 i_1417 (.A1(inputB[16]), .A2(inputA[23]), .ZN(n_1560));
   OAI21_X1 i_1419 (.A(n_1563), .B1(n_1630), .B2(n_1564), .ZN(n_1562));
   NAND2_X1 i_1420 (.A1(n_1630), .A2(n_1564), .ZN(n_1563));
   INV_X1 i_1421 (.A(n_1565), .ZN(n_1564));
   NAND2_X1 i_1422 (.A1(inputB[14]), .A2(inputA[25]), .ZN(n_1565));
   XOR2_X1 i_1423 (.A(n_1567), .B(n_1566), .Z(n_4777));
   NAND2_X1 i_1424 (.A1(inputB[13]), .A2(inputA[26]), .ZN(n_1566));
   NAND2_X1 i_1425 (.A1(n_1569), .A2(n_1568), .ZN(n_1567));
   NAND3_X1 i_1426 (.A1(inputB[11]), .A2(inputA[28]), .A3(n_1707), .ZN(n_1568));
   INV_X1 i_1427 (.A(n_1570), .ZN(n_1569));
   AOI21_X1 i_1428 (.A(n_1707), .B1(inputB[11]), .B2(inputA[28]), .ZN(n_1570));
   INV_X1 i_1429 (.A(n_1571), .ZN(n_4656));
   AOI21_X1 i_1430 (.A(n_4653), .B1(n_4652), .B2(n_1623), .ZN(n_1571));
   INV_X1 i_1431 (.A(n_1572), .ZN(n_4661));
   AOI21_X1 i_1432 (.A(n_4658), .B1(n_4657), .B2(n_1646), .ZN(n_1572));
   NOR2_X1 i_1433 (.A1(n_1653), .A2(n_1573), .ZN(n_4597));
   AOI21_X1 i_1434 (.A(n_1651), .B1(n_1811), .B2(n_1657), .ZN(n_1573));
   OAI21_X1 i_1435 (.A(n_1668), .B1(n_1672), .B2(n_1662), .ZN(n_4606));
   OAI21_X1 i_1436 (.A(n_1683), .B1(n_1687), .B2(n_1677), .ZN(n_4620));
   OAI21_X1 i_1437 (.A(n_1700), .B1(n_1702), .B2(n_1696), .ZN(n_4627));
   OAI21_X1 i_1438 (.A(n_1706), .B1(n_1709), .B2(n_1704), .ZN(n_4641));
   OAI22_X1 i_1439 (.A1(n_1853), .A2(n_1714), .B1(n_1716), .B2(n_1710), .ZN(
      n_4648));
   XOR2_X1 i_1440 (.A(n_4717), .B(n_1577), .Z(n_4719));
   XOR2_X1 i_1441 (.A(n_4707), .B(n_1582), .Z(n_1577));
   XNOR2_X1 i_1442 (.A(n_4692), .B(n_1586), .ZN(n_1582));
   INV_X1 i_1443 (.A(n_1586), .ZN(n_1583));
   AOI21_X1 i_1444 (.A(n_4531), .B1(n_4530), .B2(n_1791), .ZN(n_1586));
   INV_X1 i_1445 (.A(n_1587), .ZN(n_4589));
   AOI21_X1 i_1446 (.A(n_4586), .B1(n_4585), .B2(n_1591), .ZN(n_1587));
   INV_X1 i_1447 (.A(n_1592), .ZN(n_1591));
   AOI21_X1 i_1448 (.A(n_4436), .B1(n_4435), .B2(n_1872), .ZN(n_1592));
   XOR2_X1 i_1449 (.A(n_4712), .B(n_1597), .Z(n_4714));
   XNOR2_X1 i_1450 (.A(n_4697), .B(n_1601), .ZN(n_1597));
   INV_X1 i_1451 (.A(n_1601), .ZN(n_1598));
   AOI21_X1 i_1452 (.A(n_4556), .B1(n_4555), .B2(n_1756), .ZN(n_1601));
   INV_X1 i_1453 (.A(n_1602), .ZN(n_4579));
   AOI21_X1 i_1455 (.A(n_4576), .B1(n_4575), .B2(n_1726), .ZN(n_1602));
   XOR2_X1 i_1456 (.A(n_4702), .B(n_1607), .Z(n_4704));
   XOR2_X1 i_1457 (.A(n_4677), .B(n_1611), .Z(n_1607));
   XOR2_X1 i_1459 (.A(n_1613), .B(n_1612), .Z(n_1611));
   NAND2_X1 i_1460 (.A1(inputB[25]), .A2(inputA[13]), .ZN(n_1612));
   NAND2_X1 i_1461 (.A1(n_1616), .A2(n_1615), .ZN(n_1613));
   NAND3_X1 i_1463 (.A1(inputB[23]), .A2(inputA[15]), .A3(n_1785), .ZN(n_1615));
   INV_X1 i_1464 (.A(n_1617), .ZN(n_1616));
   AOI21_X1 i_1465 (.A(n_1785), .B1(inputB[23]), .B2(inputA[15]), .ZN(n_1617));
   INV_X1 i_1467 (.A(n_1618), .ZN(n_4574));
   AOI21_X1 i_1468 (.A(n_4571), .B1(n_4570), .B2(n_1729), .ZN(n_1618));
   INV_X1 i_1469 (.A(n_1619), .ZN(n_4569));
   AOI21_X1 i_1471 (.A(n_4566), .B1(n_4565), .B2(n_1734), .ZN(n_1619));
   XOR2_X1 i_1472 (.A(n_4687), .B(n_1622), .Z(n_4689));
   XOR2_X1 i_1473 (.A(n_4652), .B(n_1623), .Z(n_1622));
   AOI22_X1 i_1475 (.A1(n_1919), .A2(n_1839), .B1(n_1834), .B2(n_1832), .ZN(
      n_1623));
   INV_X1 i_1476 (.A(n_1624), .ZN(n_4564));
   AOI21_X1 i_1477 (.A(n_4561), .B1(n_4560), .B2(n_1727), .ZN(n_1624));
   XOR2_X1 i_1479 (.A(n_4672), .B(n_1625), .Z(n_4674));
   XOR2_X1 i_1480 (.A(n_1628), .B(n_1626), .Z(n_1625));
   NAND2_X1 i_1481 (.A1(inputB[16]), .A2(inputA[22]), .ZN(n_1626));
   NAND2_X1 i_1483 (.A1(n_1632), .A2(n_1629), .ZN(n_1628));
   NAND3_X1 i_1484 (.A1(inputB[14]), .A2(inputA[23]), .A3(n_1630), .ZN(n_1629));
   INV_X1 i_1485 (.A(n_1631), .ZN(n_1630));
   NAND2_X1 i_1486 (.A1(inputB[15]), .A2(inputA[24]), .ZN(n_1631));
   INV_X1 i_1487 (.A(n_1633), .ZN(n_1632));
   AOI22_X1 i_1488 (.A1(inputB[15]), .A2(inputA[23]), .B1(inputB[14]), .B2(
      inputA[24]), .ZN(n_1633));
   XNOR2_X1 i_1489 (.A(n_4682), .B(n_1636), .ZN(n_4684));
   INV_X1 i_1490 (.A(n_1636), .ZN(n_1634));
   AOI21_X1 i_1491 (.A(n_4526), .B1(n_4525), .B2(n_1803), .ZN(n_1636));
   INV_X1 i_1492 (.A(n_1637), .ZN(n_4554));
   AOI21_X1 i_1493 (.A(n_4551), .B1(n_4550), .B2(n_1730), .ZN(n_1637));
   XNOR2_X1 i_1494 (.A(n_4667), .B(n_1639), .ZN(n_4669));
   INV_X1 i_1495 (.A(n_1639), .ZN(n_1638));
   AOI21_X1 i_1496 (.A(n_1640), .B1(n_1798), .B2(n_1793), .ZN(n_1639));
   AOI21_X1 i_1497 (.A(n_1796), .B1(n_1797), .B2(n_1792), .ZN(n_1640));
   INV_X1 i_1498 (.A(n_1643), .ZN(n_4549));
   AOI21_X1 i_1499 (.A(n_4546), .B1(n_4545), .B2(n_1786), .ZN(n_1643));
   INV_X1 i_1500 (.A(n_1644), .ZN(n_4539));
   AOI21_X1 i_1501 (.A(n_4536), .B1(n_4535), .B2(n_1735), .ZN(n_1644));
   INV_X1 i_1502 (.A(n_1645), .ZN(n_4544));
   AOI21_X1 i_1503 (.A(n_4541), .B1(n_4540), .B2(n_1766), .ZN(n_1645));
   XOR2_X1 i_1504 (.A(n_4657), .B(n_1646), .Z(n_4659));
   OAI21_X1 i_1505 (.A(n_1822), .B1(n_1824), .B2(n_1820), .ZN(n_1646));
   XOR2_X1 i_1506 (.A(n_4662), .B(n_1649), .Z(n_4664));
   NAND2_X1 i_1507 (.A1(n_1810), .A2(n_1650), .ZN(n_1649));
   NAND2_X1 i_1508 (.A1(n_1807), .A2(n_1805), .ZN(n_1650));
   XOR2_X1 i_1509 (.A(n_1652), .B(n_1651), .Z(n_4596));
   NAND2_X1 i_1510 (.A1(inputB[31]), .A2(inputA[7]), .ZN(n_1651));
   AOI21_X1 i_1511 (.A(n_1653), .B1(n_1811), .B2(n_1657), .ZN(n_1652));
   AOI22_X1 i_1512 (.A1(inputB[30]), .A2(inputA[8]), .B1(inputB[29]), .B2(
      inputA[9]), .ZN(n_1653));
   INV_X1 i_1513 (.A(n_1658), .ZN(n_1657));
   NAND2_X1 i_1514 (.A1(inputB[30]), .A2(inputA[9]), .ZN(n_1658));
   XOR2_X1 i_1515 (.A(n_1667), .B(n_1662), .Z(n_4605));
   NAND2_X1 i_1516 (.A1(inputB[28]), .A2(inputA[10]), .ZN(n_1662));
   NAND2_X1 i_1517 (.A1(n_1671), .A2(n_1668), .ZN(n_1667));
   NAND4_X1 i_1518 (.A1(inputB[26]), .A2(inputA[11]), .A3(inputB[27]), .A4(
      inputA[12]), .ZN(n_1668));
   INV_X1 i_1519 (.A(n_1672), .ZN(n_1671));
   AOI22_X1 i_1520 (.A1(inputB[27]), .A2(inputA[11]), .B1(inputB[26]), .B2(
      inputA[12]), .ZN(n_1672));
   XOR2_X1 i_1521 (.A(n_1682), .B(n_1677), .Z(n_4619));
   NAND2_X1 i_1522 (.A1(inputB[22]), .A2(inputA[16]), .ZN(n_1677));
   NAND2_X1 i_1523 (.A1(n_1686), .A2(n_1683), .ZN(n_1682));
   NAND3_X1 i_1524 (.A1(inputB[21]), .A2(inputA[17]), .A3(n_1692), .ZN(n_1683));
   INV_X1 i_1525 (.A(n_1687), .ZN(n_1686));
   AOI21_X1 i_1527 (.A(n_1692), .B1(inputB[21]), .B2(inputA[17]), .ZN(n_1687));
   AND2_X1 i_1528 (.A1(inputB[20]), .A2(inputA[18]), .ZN(n_1692));
   XOR2_X1 i_1529 (.A(n_1697), .B(n_1696), .Z(n_4626));
   NAND2_X1 i_1531 (.A1(inputB[19]), .A2(inputA[19]), .ZN(n_1696));
   NAND2_X1 i_1532 (.A1(n_1701), .A2(n_1700), .ZN(n_1697));
   NAND3_X1 i_1533 (.A1(inputB[18]), .A2(inputA[20]), .A3(n_1703), .ZN(n_1700));
   INV_X1 i_1535 (.A(n_1702), .ZN(n_1701));
   AOI21_X1 i_1536 (.A(n_1703), .B1(inputB[18]), .B2(inputA[20]), .ZN(n_1702));
   AND2_X1 i_1537 (.A1(inputB[17]), .A2(inputA[21]), .ZN(n_1703));
   XOR2_X1 i_1539 (.A(n_1705), .B(n_1704), .Z(n_4640));
   NAND2_X1 i_1540 (.A1(inputB[13]), .A2(inputA[25]), .ZN(n_1704));
   NAND2_X1 i_1541 (.A1(n_1708), .A2(n_1706), .ZN(n_1705));
   NAND2_X1 i_1543 (.A1(n_1838), .A2(n_1707), .ZN(n_1706));
   AND2_X1 i_1544 (.A1(inputB[12]), .A2(inputA[27]), .ZN(n_1707));
   INV_X1 i_1545 (.A(n_1709), .ZN(n_1708));
   AOI22_X1 i_1547 (.A1(inputB[12]), .A2(inputA[26]), .B1(inputB[11]), .B2(
      inputA[27]), .ZN(n_1709));
   XOR2_X1 i_1548 (.A(n_1711), .B(n_1710), .Z(n_4647));
   NAND2_X1 i_1549 (.A1(inputB[10]), .A2(inputA[28]), .ZN(n_1710));
   OAI21_X1 i_1551 (.A(n_1715), .B1(n_1853), .B2(n_1714), .ZN(n_1711));
   NAND2_X1 i_1552 (.A1(inputB[9]), .A2(inputA[30]), .ZN(n_1714));
   INV_X1 i_1553 (.A(n_1716), .ZN(n_1715));
   AOI22_X1 i_1555 (.A1(inputB[9]), .A2(inputA[29]), .B1(inputB[8]), .B2(
      inputA[30]), .ZN(n_1716));
   INV_X1 i_1556 (.A(n_1717), .ZN(n_4519));
   AOI21_X1 i_1557 (.A(n_4516), .B1(n_4515), .B2(n_1731), .ZN(n_1717));
   INV_X1 i_1558 (.A(n_1718), .ZN(n_4524));
   AOI21_X1 i_1559 (.A(n_4521), .B1(n_4520), .B2(n_1801), .ZN(n_1718));
   OAI21_X1 i_1560 (.A(n_1817), .B1(n_1819), .B2(n_1813), .ZN(n_4461));
   OAI21_X1 i_1561 (.A(n_1781), .B1(n_1776), .B2(n_1767), .ZN(n_4468));
   OAI21_X1 i_1562 (.A(n_1827), .B1(n_1831), .B2(n_1825), .ZN(n_4482));
   OAI21_X1 i_1563 (.A(n_1741), .B1(n_1746), .B2(n_1745), .ZN(n_4489));
   AOI22_X1 i_1564 (.A1(n_2003), .A2(n_1853), .B1(n_1847), .B2(n_1843), .ZN(
      n_4503));
   NAND2_X1 i_1565 (.A1(inputB[7]), .A2(inputA[31]), .ZN(n_383));
   XNOR2_X1 i_1566 (.A(n_4580), .B(n_1722), .ZN(n_4582));
   INV_X1 i_1567 (.A(n_1722), .ZN(n_1721));
   AOI21_X1 i_1568 (.A(n_4431), .B1(n_4430), .B2(n_1882), .ZN(n_1722));
   INV_X1 i_1569 (.A(n_1723), .ZN(n_4444));
   AOI21_X1 i_1570 (.A(n_4441), .B1(n_4440), .B2(n_1724), .ZN(n_1723));
   INV_X1 i_1571 (.A(n_1725), .ZN(n_1724));
   AOI21_X1 i_1572 (.A(n_4286), .B1(n_4285), .B2(n_2019), .ZN(n_1725));
   XOR2_X1 i_1573 (.A(n_4575), .B(n_1726), .Z(n_4577));
   XNOR2_X1 i_1574 (.A(n_4560), .B(n_1728), .ZN(n_1726));
   INV_X1 i_1575 (.A(n_1728), .ZN(n_1727));
   AOI21_X1 i_1576 (.A(n_4401), .B1(n_4400), .B2(n_1906), .ZN(n_1728));
   XOR2_X1 i_1577 (.A(n_4570), .B(n_1729), .Z(n_4572));
   XOR2_X1 i_1578 (.A(n_4550), .B(n_1730), .Z(n_1729));
   XOR2_X1 i_1579 (.A(n_4515), .B(n_1731), .Z(n_1730));
   AOI21_X1 i_1580 (.A(n_1732), .B1(n_2056), .B2(n_1997), .ZN(n_1731));
   NOR2_X1 i_1581 (.A1(n_1996), .A2(n_1992), .ZN(n_1732));
   XOR2_X1 i_1582 (.A(n_4565), .B(n_1734), .Z(n_4567));
   XOR2_X1 i_1583 (.A(n_4535), .B(n_1735), .Z(n_1734));
   XNOR2_X1 i_1584 (.A(n_1746), .B(n_1736), .ZN(n_1735));
   NOR2_X1 i_1585 (.A1(n_1745), .A2(n_1737), .ZN(n_1736));
   INV_X1 i_1586 (.A(n_1741), .ZN(n_1737));
   NAND4_X1 i_1587 (.A1(inputB[14]), .A2(inputA[22]), .A3(inputB[15]), .A4(
      inputA[23]), .ZN(n_1741));
   AOI22_X1 i_1588 (.A1(inputB[15]), .A2(inputA[22]), .B1(inputB[14]), .B2(
      inputA[23]), .ZN(n_1745));
   NAND2_X1 i_1589 (.A1(inputB[16]), .A2(inputA[21]), .ZN(n_1746));
   INV_X1 i_1590 (.A(n_1747), .ZN(n_4429));
   AOI21_X1 i_1591 (.A(n_4426), .B1(n_4425), .B2(n_1893), .ZN(n_1747));
   INV_X1 i_1592 (.A(n_1750), .ZN(n_4424));
   AOI21_X1 i_1593 (.A(n_4421), .B1(n_4420), .B2(n_1895), .ZN(n_1750));
   INV_X1 i_1594 (.A(n_1751), .ZN(n_4419));
   AOI21_X1 i_1595 (.A(n_4416), .B1(n_4415), .B2(n_1883), .ZN(n_1751));
   XNOR2_X1 i_1596 (.A(n_4555), .B(n_1757), .ZN(n_4557));
   INV_X1 i_1597 (.A(n_1757), .ZN(n_1756));
   AOI21_X1 i_1599 (.A(n_4386), .B1(n_4385), .B2(n_1910), .ZN(n_1757));
   INV_X1 i_1600 (.A(n_1761), .ZN(n_4414));
   AOI21_X1 i_1601 (.A(n_4411), .B1(n_4410), .B2(n_1902), .ZN(n_1761));
   XOR2_X1 i_1603 (.A(n_4540), .B(n_1766), .Z(n_4542));
   XOR2_X1 i_1604 (.A(n_1771), .B(n_1767), .Z(n_1766));
   NAND2_X1 i_1605 (.A1(inputB[25]), .A2(inputA[12]), .ZN(n_1767));
   NAND2_X1 i_1607 (.A1(n_1781), .A2(n_1775), .ZN(n_1771));
   INV_X1 i_1608 (.A(n_1776), .ZN(n_1775));
   AOI22_X1 i_1609 (.A1(inputB[24]), .A2(inputA[13]), .B1(inputB[23]), .B2(
      inputA[14]), .ZN(n_1776));
   NAND3_X1 i_1611 (.A1(inputB[23]), .A2(inputA[13]), .A3(n_1785), .ZN(n_1781));
   AND2_X1 i_1612 (.A1(inputB[24]), .A2(inputA[14]), .ZN(n_1785));
   XNOR2_X1 i_1613 (.A(n_4545), .B(n_1789), .ZN(n_4547));
   INV_X1 i_1615 (.A(n_1789), .ZN(n_1786));
   AOI21_X1 i_1616 (.A(n_4381), .B1(n_4380), .B2(n_1903), .ZN(n_1789));
   INV_X1 i_1617 (.A(n_1790), .ZN(n_4409));
   AOI21_X1 i_1619 (.A(n_4406), .B1(n_4405), .B2(n_1908), .ZN(n_1790));
   XOR2_X1 i_1620 (.A(n_4530), .B(n_1791), .Z(n_4532));
   XOR2_X1 i_1621 (.A(n_1798), .B(n_1792), .Z(n_1791));
   XNOR2_X1 i_1623 (.A(n_1796), .B(n_1793), .ZN(n_1792));
   NAND2_X1 i_1624 (.A1(inputB[6]), .A2(inputA[31]), .ZN(n_1793));
   NAND2_X1 i_1625 (.A1(inputB[7]), .A2(inputA[30]), .ZN(n_1796));
   INV_X1 i_1627 (.A(n_1798), .ZN(n_1797));
   AOI21_X1 i_1628 (.A(n_2009), .B1(n_2010), .B2(n_2006), .ZN(n_1798));
   INV_X1 i_1629 (.A(n_1799), .ZN(n_4394));
   AOI21_X1 i_1631 (.A(n_4391), .B1(n_4390), .B2(n_1921), .ZN(n_1799));
   INV_X1 i_1632 (.A(n_1800), .ZN(n_4399));
   AOI21_X1 i_1633 (.A(n_4396), .B1(n_4395), .B2(n_1885), .ZN(n_1800));
   XOR2_X1 i_1634 (.A(n_4520), .B(n_1801), .Z(n_4522));
   AOI21_X1 i_1635 (.A(n_1802), .B1(n_2070), .B2(n_1985), .ZN(n_1801));
   NOR2_X1 i_1636 (.A1(n_1984), .A2(n_1975), .ZN(n_1802));
   XNOR2_X1 i_1637 (.A(n_4525), .B(n_1804), .ZN(n_4527));
   INV_X1 i_1638 (.A(n_1804), .ZN(n_1803));
   AOI21_X1 i_1639 (.A(n_4376), .B1(n_4375), .B2(n_1950), .ZN(n_1804));
   XOR2_X1 i_1640 (.A(n_1806), .B(n_1805), .Z(n_4451));
   NAND2_X1 i_1641 (.A1(inputB[31]), .A2(inputA[6]), .ZN(n_1805));
   AND2_X1 i_1642 (.A1(n_1810), .A2(n_1807), .ZN(n_1806));
   NAND2_X1 i_1643 (.A1(n_1890), .A2(n_1812), .ZN(n_1807));
   NAND2_X1 i_1644 (.A1(n_1889), .A2(n_1811), .ZN(n_1810));
   INV_X1 i_1645 (.A(n_1812), .ZN(n_1811));
   NAND2_X1 i_1646 (.A1(inputB[29]), .A2(inputA[8]), .ZN(n_1812));
   XOR2_X1 i_1647 (.A(n_1814), .B(n_1813), .Z(n_4460));
   NAND2_X1 i_1648 (.A1(inputB[28]), .A2(inputA[9]), .ZN(n_1813));
   NAND2_X1 i_1649 (.A1(n_1818), .A2(n_1817), .ZN(n_1814));
   NAND4_X1 i_1650 (.A1(inputB[26]), .A2(inputA[10]), .A3(inputB[27]), .A4(
      inputA[11]), .ZN(n_1817));
   INV_X1 i_1651 (.A(n_1819), .ZN(n_1818));
   AOI22_X1 i_1652 (.A1(inputB[27]), .A2(inputA[10]), .B1(inputB[26]), .B2(
      inputA[11]), .ZN(n_1819));
   XOR2_X1 i_1653 (.A(n_1821), .B(n_1820), .Z(n_4474));
   NAND2_X1 i_1654 (.A1(inputB[22]), .A2(inputA[15]), .ZN(n_1820));
   NAND2_X1 i_1655 (.A1(n_1823), .A2(n_1822), .ZN(n_1821));
   NAND3_X1 i_1656 (.A1(inputB[20]), .A2(inputA[17]), .A3(n_1929), .ZN(n_1822));
   INV_X1 i_1657 (.A(n_1824), .ZN(n_1823));
   AOI21_X1 i_1658 (.A(n_1929), .B1(inputB[20]), .B2(inputA[17]), .ZN(n_1824));
   XOR2_X1 i_1659 (.A(n_1826), .B(n_1825), .Z(n_4481));
   NAND2_X1 i_1660 (.A1(inputB[19]), .A2(inputA[18]), .ZN(n_1825));
   NAND2_X1 i_1661 (.A1(n_1828), .A2(n_1827), .ZN(n_1826));
   NAND4_X1 i_1662 (.A1(inputB[18]), .A2(inputA[19]), .A3(inputB[17]), .A4(
      inputA[20]), .ZN(n_1827));
   INV_X1 i_1663 (.A(n_1831), .ZN(n_1828));
   AOI22_X1 i_1664 (.A1(inputB[18]), .A2(inputA[19]), .B1(inputB[17]), .B2(
      inputA[20]), .ZN(n_1831));
   XOR2_X1 i_1665 (.A(n_1833), .B(n_1832), .Z(n_4495));
   NAND2_X1 i_1666 (.A1(inputB[13]), .A2(inputA[24]), .ZN(n_1832));
   OAI21_X1 i_1667 (.A(n_1834), .B1(n_1918), .B2(n_1838), .ZN(n_1833));
   NAND2_X1 i_1668 (.A1(n_1918), .A2(n_1838), .ZN(n_1834));
   INV_X1 i_1669 (.A(n_1839), .ZN(n_1838));
   NAND2_X1 i_1670 (.A1(inputB[11]), .A2(inputA[26]), .ZN(n_1839));
   XOR2_X1 i_1671 (.A(n_1844), .B(n_1843), .Z(n_4502));
   NAND2_X1 i_1672 (.A1(inputB[10]), .A2(inputA[27]), .ZN(n_1843));
   OAI21_X1 i_1674 (.A(n_1847), .B1(n_2002), .B2(n_1848), .ZN(n_1844));
   NAND2_X1 i_1675 (.A1(n_2002), .A2(n_1848), .ZN(n_1847));
   INV_X1 i_1676 (.A(n_1853), .ZN(n_1848));
   NAND2_X1 i_1678 (.A1(inputB[8]), .A2(inputA[29]), .ZN(n_1853));
   INV_X1 i_1679 (.A(n_1858), .ZN(n_4369));
   AOI21_X1 i_1680 (.A(n_4366), .B1(n_4365), .B2(n_1945), .ZN(n_1858));
   INV_X1 i_1682 (.A(n_1862), .ZN(n_4374));
   AOI21_X1 i_1683 (.A(n_4371), .B1(n_4370), .B2(n_1907), .ZN(n_1862));
   INV_X1 i_1684 (.A(n_1863), .ZN(n_4302));
   AOI22_X1 i_1686 (.A1(n_2108), .A2(n_1889), .B1(n_1887), .B2(n_1886), .ZN(
      n_1863));
   OAI21_X1 i_1687 (.A(n_1965), .B1(n_1974), .B2(n_1960), .ZN(n_4311));
   OAI21_X1 i_1688 (.A(n_1928), .B1(n_1927), .B2(n_1922), .ZN(n_4325));
   OAI21_X1 i_1690 (.A(n_1989), .B1(n_1991), .B2(n_1986), .ZN(n_4332));
   OAI21_X1 i_1691 (.A(n_1917), .B1(n_1916), .B2(n_1911), .ZN(n_4346));
   OAI21_X1 i_1692 (.A(n_2001), .B1(n_2005), .B2(n_1998), .ZN(n_4353));
   INV_X1 i_1694 (.A(n_1864), .ZN(n_4294));
   AOI21_X1 i_1695 (.A(n_4291), .B1(n_4290), .B2(n_1868), .ZN(n_1864));
   XOR2_X1 i_1696 (.A(n_4280), .B(n_1878), .Z(n_1868));
   XNOR2_X1 i_1698 (.A(n_4435), .B(n_1873), .ZN(n_4437));
   INV_X1 i_1699 (.A(n_1873), .ZN(n_1872));
   AOI21_X1 i_1700 (.A(n_4281), .B1(n_4280), .B2(n_1878), .ZN(n_1873));
   XNOR2_X1 i_1702 (.A(n_4260), .B(n_1898), .ZN(n_1878));
   XOR2_X1 i_1703 (.A(n_4430), .B(n_1882), .Z(n_4432));
   XOR2_X1 i_1704 (.A(n_4415), .B(n_1883), .Z(n_1882));
   XOR2_X1 i_1706 (.A(n_4395), .B(n_1885), .Z(n_1883));
   XOR2_X1 i_1707 (.A(n_1887), .B(n_1886), .Z(n_1885));
   NAND2_X1 i_1708 (.A1(inputB[31]), .A2(inputA[5]), .ZN(n_1886));
   AOI21_X1 i_1710 (.A(n_1888), .B1(n_2108), .B2(n_1889), .ZN(n_1887));
   AOI22_X1 i_1711 (.A1(inputB[30]), .A2(inputA[6]), .B1(inputB[29]), .B2(
      inputA[7]), .ZN(n_1888));
   INV_X1 i_1712 (.A(n_1890), .ZN(n_1889));
   NAND2_X1 i_1713 (.A1(inputB[30]), .A2(inputA[7]), .ZN(n_1890));
   XNOR2_X1 i_1714 (.A(n_4425), .B(n_1894), .ZN(n_4427));
   INV_X1 i_1715 (.A(n_1894), .ZN(n_1893));
   AOI21_X1 i_1716 (.A(n_4266), .B1(n_4265), .B2(n_2028), .ZN(n_1894));
   XNOR2_X1 i_1717 (.A(n_4420), .B(n_1896), .ZN(n_4422));
   INV_X1 i_1718 (.A(n_1896), .ZN(n_1895));
   AOI21_X1 i_1719 (.A(n_4261), .B1(n_4260), .B2(n_1897), .ZN(n_1896));
   INV_X1 i_1720 (.A(n_1898), .ZN(n_1897));
   AOI21_X1 i_1721 (.A(n_4102), .B1(n_4101), .B2(n_2210), .ZN(n_1898));
   INV_X1 i_1722 (.A(n_1900), .ZN(n_4279));
   AOI21_X1 i_1723 (.A(n_4276), .B1(n_4275), .B2(n_2023), .ZN(n_1900));
   INV_X1 i_1724 (.A(n_1901), .ZN(n_4274));
   AOI21_X1 i_1725 (.A(n_4271), .B1(n_4270), .B2(n_2025), .ZN(n_1901));
   XOR2_X1 i_1726 (.A(n_4410), .B(n_1902), .Z(n_4412));
   XNOR2_X1 i_1727 (.A(n_4380), .B(n_1904), .ZN(n_1902));
   INV_X1 i_1728 (.A(n_1904), .ZN(n_1903));
   AOI21_X1 i_1729 (.A(n_4211), .B1(n_4210), .B2(n_2035), .ZN(n_1904));
   XOR2_X1 i_1730 (.A(n_4400), .B(n_1906), .Z(n_4402));
   XOR2_X1 i_1731 (.A(n_4370), .B(n_1907), .Z(n_1906));
   OAI21_X1 i_1732 (.A(n_2118), .B1(n_2122), .B2(n_2116), .ZN(n_1907));
   XNOR2_X1 i_1733 (.A(n_4405), .B(n_1909), .ZN(n_4407));
   INV_X1 i_1734 (.A(n_1909), .ZN(n_1908));
   AOI21_X1 i_1735 (.A(n_4236), .B1(n_4235), .B2(n_2042), .ZN(n_1909));
   XOR2_X1 i_1736 (.A(n_4385), .B(n_1910), .Z(n_4387));
   XOR2_X1 i_1737 (.A(n_1914), .B(n_1911), .Z(n_1910));
   NAND2_X1 i_1738 (.A1(inputB[13]), .A2(inputA[23]), .ZN(n_1911));
   NAND2_X1 i_1739 (.A1(n_1917), .A2(n_1915), .ZN(n_1914));
   INV_X1 i_1740 (.A(n_1916), .ZN(n_1915));
   AOI22_X1 i_1741 (.A1(inputB[12]), .A2(inputA[24]), .B1(inputB[11]), .B2(
      inputA[25]), .ZN(n_1916));
   NAND2_X1 i_1742 (.A1(n_2136), .A2(n_1918), .ZN(n_1917));
   INV_X1 i_1743 (.A(n_1919), .ZN(n_1918));
   NAND2_X1 i_1744 (.A1(inputB[12]), .A2(inputA[25]), .ZN(n_1919));
   XOR2_X1 i_1745 (.A(n_4390), .B(n_1921), .Z(n_4392));
   XOR2_X1 i_1746 (.A(n_1923), .B(n_1922), .Z(n_1921));
   NAND2_X1 i_1747 (.A1(inputB[22]), .A2(inputA[14]), .ZN(n_1922));
   NAND2_X1 i_1748 (.A1(n_1928), .A2(n_1924), .ZN(n_1923));
   INV_X1 i_1749 (.A(n_1927), .ZN(n_1924));
   AOI22_X1 i_1750 (.A1(inputB[21]), .A2(inputA[15]), .B1(inputB[20]), .B2(
      inputA[16]), .ZN(n_1927));
   NAND2_X1 i_1751 (.A1(n_2123), .A2(n_1929), .ZN(n_1928));
   AND2_X1 i_1752 (.A1(inputB[21]), .A2(inputA[16]), .ZN(n_1929));
   INV_X1 i_1753 (.A(n_1930), .ZN(n_4254));
   AOI21_X1 i_1754 (.A(n_4251), .B1(n_4250), .B2(n_2032), .ZN(n_1930));
   INV_X1 i_1755 (.A(n_1931), .ZN(n_4259));
   AOI21_X1 i_1756 (.A(n_4256), .B1(n_4255), .B2(n_2036), .ZN(n_1931));
   INV_X1 i_1757 (.A(n_1935), .ZN(n_4249));
   AOI21_X1 i_1758 (.A(n_4246), .B1(n_4245), .B2(n_2029), .ZN(n_1935));
   INV_X1 i_1759 (.A(n_1939), .ZN(n_4234));
   AOI21_X1 i_1761 (.A(n_4231), .B1(n_4230), .B2(n_2086), .ZN(n_1939));
   INV_X1 i_1762 (.A(n_1940), .ZN(n_4244));
   AOI21_X1 i_1763 (.A(n_4241), .B1(n_4240), .B2(n_2057), .ZN(n_1940));
   XOR2_X1 i_1765 (.A(n_4365), .B(n_1945), .Z(n_4367));
   OAI21_X1 i_1766 (.A(n_2132), .B1(n_2135), .B2(n_2130), .ZN(n_1945));
   XOR2_X1 i_1767 (.A(n_4375), .B(n_1950), .Z(n_4377));
   NAND2_X1 i_1769 (.A1(n_2106), .A2(n_1954), .ZN(n_1950));
   NAND2_X1 i_1770 (.A1(n_2105), .A2(n_2103), .ZN(n_1954));
   INV_X1 i_1771 (.A(n_1955), .ZN(n_4229));
   AOI21_X1 i_1773 (.A(n_4226), .B1(n_4225), .B2(n_2080), .ZN(n_1955));
   XOR2_X1 i_1774 (.A(n_1964), .B(n_1960), .Z(n_4310));
   NAND2_X1 i_1775 (.A1(inputB[28]), .A2(inputA[8]), .ZN(n_1960));
   NAND2_X1 i_1777 (.A1(n_1970), .A2(n_1965), .ZN(n_1964));
   NAND3_X1 i_1778 (.A1(inputB[27]), .A2(inputA[10]), .A3(n_2114), .ZN(n_1965));
   INV_X1 i_1779 (.A(n_1974), .ZN(n_1970));
   AOI22_X1 i_1781 (.A1(inputB[27]), .A2(inputA[9]), .B1(inputB[26]), .B2(
      inputA[10]), .ZN(n_1974));
   XOR2_X1 i_1782 (.A(n_1980), .B(n_1975), .Z(n_4317));
   AND2_X1 i_1783 (.A1(inputB[25]), .A2(inputA[11]), .ZN(n_1975));
   AOI21_X1 i_1785 (.A(n_1984), .B1(n_2070), .B2(n_1985), .ZN(n_1980));
   NOR2_X1 i_1786 (.A1(n_2070), .A2(n_1985), .ZN(n_1984));
   NAND2_X1 i_1787 (.A1(inputB[23]), .A2(inputA[13]), .ZN(n_1985));
   XOR2_X1 i_1789 (.A(n_1988), .B(n_1986), .Z(n_4331));
   NAND2_X1 i_1790 (.A1(inputB[19]), .A2(inputA[17]), .ZN(n_1986));
   NAND2_X1 i_1791 (.A1(n_1990), .A2(n_1989), .ZN(n_1988));
   NAND4_X1 i_1793 (.A1(inputB[18]), .A2(inputA[18]), .A3(inputB[17]), .A4(
      inputA[19]), .ZN(n_1989));
   INV_X1 i_1794 (.A(n_1991), .ZN(n_1990));
   AOI22_X1 i_1795 (.A1(inputB[18]), .A2(inputA[18]), .B1(inputB[17]), .B2(
      inputA[19]), .ZN(n_1991));
   XOR2_X1 i_1797 (.A(n_1995), .B(n_1992), .Z(n_4338));
   AND2_X1 i_1798 (.A1(inputB[16]), .A2(inputA[20]), .ZN(n_1992));
   AOI21_X1 i_1799 (.A(n_1996), .B1(n_2056), .B2(n_1997), .ZN(n_1995));
   NOR2_X1 i_1800 (.A1(n_2056), .A2(n_1997), .ZN(n_1996));
   NAND2_X1 i_1801 (.A1(inputB[14]), .A2(inputA[22]), .ZN(n_1997));
   XOR2_X1 i_1802 (.A(n_1999), .B(n_1998), .Z(n_4352));
   NAND2_X1 i_1803 (.A1(inputB[10]), .A2(inputA[26]), .ZN(n_1998));
   NAND2_X1 i_1804 (.A1(n_2004), .A2(n_2001), .ZN(n_1999));
   NAND3_X1 i_1805 (.A1(inputB[8]), .A2(inputA[27]), .A3(n_2002), .ZN(n_2001));
   INV_X1 i_1806 (.A(n_2003), .ZN(n_2002));
   NAND2_X1 i_1807 (.A1(inputB[9]), .A2(inputA[28]), .ZN(n_2003));
   INV_X1 i_1808 (.A(n_2005), .ZN(n_2004));
   AOI22_X1 i_1809 (.A1(inputB[9]), .A2(inputA[27]), .B1(inputB[8]), .B2(
      inputA[28]), .ZN(n_2005));
   XNOR2_X1 i_1810 (.A(n_2007), .B(n_2006), .ZN(n_4358));
   NAND2_X1 i_1811 (.A1(inputB[7]), .A2(inputA[29]), .ZN(n_2006));
   NOR2_X1 i_1812 (.A1(n_2011), .A2(n_2009), .ZN(n_2007));
   AND3_X1 i_1813 (.A1(inputB[5]), .A2(inputA[31]), .A3(n_2096), .ZN(n_2009));
   INV_X1 i_1814 (.A(n_2011), .ZN(n_2010));
   AOI21_X1 i_1815 (.A(n_2096), .B1(inputB[5]), .B2(inputA[31]), .ZN(n_2011));
   INV_X1 i_1816 (.A(n_2012), .ZN(n_4219));
   AOI21_X1 i_1817 (.A(n_4216), .B1(n_4215), .B2(n_2101), .ZN(n_2012));
   INV_X1 i_1818 (.A(n_2013), .ZN(n_4224));
   AOI21_X1 i_1819 (.A(n_4221), .B1(n_4220), .B2(n_2102), .ZN(n_2013));
   AOI22_X1 i_1820 (.A1(n_2233), .A2(n_2115), .B1(n_2112), .B2(n_2110), .ZN(
      n_4157));
   OAI22_X1 i_1821 (.A1(n_2258), .A2(n_2070), .B1(n_2066), .B2(n_2060), .ZN(
      n_4164));
   OAI21_X1 i_1822 (.A(n_2126), .B1(n_2129), .B2(n_2124), .ZN(n_4178));
   OAI22_X1 i_1823 (.A1(n_2284), .A2(n_2056), .B1(n_2055), .B2(n_2045), .ZN(
      n_4185));
   OAI21_X1 i_1824 (.A(n_2139), .B1(n_2143), .B2(n_2137), .ZN(n_4199));
   AOI21_X1 i_1825 (.A(n_2094), .B1(n_2095), .B2(n_2090), .ZN(n_4206));
   INV_X1 i_1826 (.A(n_2016), .ZN(n_4140));
   AOI21_X1 i_1827 (.A(n_4137), .B1(n_4136), .B2(n_2017), .ZN(n_2016));
   INV_X1 i_1828 (.A(n_2018), .ZN(n_2017));
   AOI21_X1 i_1829 (.A(n_3970), .B1(n_3969), .B2(n_2334), .ZN(n_2018));
   XNOR2_X1 i_1830 (.A(n_4285), .B(n_2020), .ZN(n_4287));
   INV_X1 i_1831 (.A(n_2020), .ZN(n_2019));
   AOI21_X1 i_1832 (.A(n_4127), .B1(n_4126), .B2(n_2161), .ZN(n_2020));
   INV_X1 i_1833 (.A(n_2022), .ZN(n_4135));
   AOI21_X1 i_1834 (.A(n_4132), .B1(n_4131), .B2(n_2159), .ZN(n_2022));
   XNOR2_X1 i_1835 (.A(n_4275), .B(n_2024), .ZN(n_4277));
   INV_X1 i_1836 (.A(n_2024), .ZN(n_2023));
   AOI21_X1 i_1837 (.A(n_4112), .B1(n_4111), .B2(n_2180), .ZN(n_2024));
   XNOR2_X1 i_1838 (.A(n_4270), .B(n_2026), .ZN(n_4272));
   INV_X1 i_1839 (.A(n_2026), .ZN(n_2025));
   AOI21_X1 i_1840 (.A(n_4107), .B1(n_4106), .B2(n_2204), .ZN(n_2026));
   INV_X1 i_1841 (.A(n_2027), .ZN(n_4125));
   AOI21_X1 i_1842 (.A(n_4122), .B1(n_4121), .B2(n_2170), .ZN(n_2027));
   XOR2_X1 i_1843 (.A(n_4265), .B(n_2028), .Z(n_4267));
   XNOR2_X1 i_1844 (.A(n_4245), .B(n_2030), .ZN(n_2028));
   INV_X1 i_1845 (.A(n_2030), .ZN(n_2029));
   AOI21_X1 i_1846 (.A(n_4072), .B1(n_4071), .B2(n_2235), .ZN(n_2030));
   INV_X1 i_1848 (.A(n_2031), .ZN(n_4120));
   AOI21_X1 i_1849 (.A(n_4117), .B1(n_4116), .B2(n_2174), .ZN(n_2031));
   XOR2_X1 i_1850 (.A(n_4250), .B(n_2032), .Z(n_4252));
   XOR2_X1 i_1852 (.A(n_4210), .B(n_2035), .Z(n_2032));
   OAI22_X1 i_1853 (.A1(n_2460), .A2(n_2195), .B1(n_2190), .B2(n_2185), .ZN(
      n_2035));
   XNOR2_X1 i_1854 (.A(n_4255), .B(n_2041), .ZN(n_4257));
   INV_X1 i_1856 (.A(n_2041), .ZN(n_2036));
   AOI21_X1 i_1857 (.A(n_4077), .B1(n_4076), .B2(n_2184), .ZN(n_2041));
   XOR2_X1 i_1858 (.A(n_4235), .B(n_2042), .Z(n_4237));
   XOR2_X1 i_1860 (.A(n_2046), .B(n_2045), .Z(n_2042));
   NAND2_X1 i_1861 (.A1(inputB[16]), .A2(inputA[19]), .ZN(n_2045));
   OAI21_X1 i_1862 (.A(n_2051), .B1(n_2284), .B2(n_2056), .ZN(n_2046));
   INV_X1 i_1864 (.A(n_2055), .ZN(n_2051));
   AOI22_X1 i_1865 (.A1(inputB[15]), .A2(inputA[20]), .B1(inputB[14]), .B2(
      inputA[21]), .ZN(n_2055));
   NAND2_X1 i_1866 (.A1(inputB[15]), .A2(inputA[21]), .ZN(n_2056));
   XOR2_X1 i_1868 (.A(n_4240), .B(n_2057), .Z(n_4242));
   XOR2_X1 i_1869 (.A(n_2061), .B(n_2060), .Z(n_2057));
   NAND2_X1 i_1870 (.A1(inputB[25]), .A2(inputA[10]), .ZN(n_2060));
   OAI21_X1 i_1872 (.A(n_2062), .B1(n_2258), .B2(n_2070), .ZN(n_2061));
   INV_X1 i_1873 (.A(n_2066), .ZN(n_2062));
   AOI22_X1 i_1874 (.A1(inputB[24]), .A2(inputA[11]), .B1(inputB[23]), .B2(
      inputA[12]), .ZN(n_2066));
   NAND2_X1 i_1876 (.A1(inputB[24]), .A2(inputA[12]), .ZN(n_2070));
   INV_X1 i_1877 (.A(n_2071), .ZN(n_4095));
   AOI21_X1 i_1878 (.A(n_4092), .B1(n_4091), .B2(n_2213), .ZN(n_2071));
   INV_X1 i_1880 (.A(n_2076), .ZN(n_4100));
   AOI21_X1 i_1881 (.A(n_4097), .B1(n_4096), .B2(n_2208), .ZN(n_2076));
   XNOR2_X1 i_1882 (.A(n_4225), .B(n_2081), .ZN(n_4227));
   INV_X1 i_1884 (.A(n_2081), .ZN(n_2080));
   AOI21_X1 i_1885 (.A(n_4062), .B1(n_4061), .B2(n_2240), .ZN(n_2081));
   XOR2_X1 i_1886 (.A(n_4230), .B(n_2086), .Z(n_4232));
   XOR2_X1 i_1888 (.A(n_2091), .B(n_2090), .Z(n_2086));
   NAND2_X1 i_1889 (.A1(inputB[7]), .A2(inputA[28]), .ZN(n_2090));
   NAND2_X1 i_1890 (.A1(n_2095), .A2(n_2093), .ZN(n_2091));
   INV_X1 i_1891 (.A(n_2094), .ZN(n_2093));
   AOI22_X1 i_1892 (.A1(inputB[6]), .A2(inputA[29]), .B1(inputB[5]), .B2(
      inputA[30]), .ZN(n_2094));
   OR2_X1 i_1893 (.A1(n_2309), .A2(n_2096), .ZN(n_2095));
   NAND2_X1 i_1894 (.A1(inputB[6]), .A2(inputA[30]), .ZN(n_2096));
   INV_X1 i_1895 (.A(n_2097), .ZN(n_4085));
   AOI21_X1 i_1896 (.A(n_4082), .B1(n_4081), .B2(n_2215), .ZN(n_2097));
   INV_X1 i_1897 (.A(n_2098), .ZN(n_4090));
   AOI21_X1 i_1898 (.A(n_4087), .B1(n_4086), .B2(n_2224), .ZN(n_2098));
   XOR2_X1 i_1899 (.A(n_4215), .B(n_2101), .Z(n_4217));
   AOI21_X1 i_1900 (.A(n_2219), .B1(n_2222), .B2(n_2216), .ZN(n_2101));
   XOR2_X1 i_1901 (.A(n_4220), .B(n_2102), .Z(n_4222));
   AOI21_X1 i_1902 (.A(n_2230), .B1(n_2231), .B2(n_2225), .ZN(n_2102));
   XOR2_X1 i_1903 (.A(n_2104), .B(n_2103), .Z(n_4147));
   NAND2_X1 i_1904 (.A1(inputB[31]), .A2(inputA[4]), .ZN(n_2103));
   AND2_X1 i_1905 (.A1(n_2106), .A2(n_2105), .ZN(n_2104));
   NAND2_X1 i_1906 (.A1(n_2247), .A2(n_2109), .ZN(n_2105));
   NAND2_X1 i_1907 (.A1(n_2246), .A2(n_2108), .ZN(n_2106));
   INV_X1 i_1908 (.A(n_2109), .ZN(n_2108));
   NAND2_X1 i_1909 (.A1(inputB[29]), .A2(inputA[6]), .ZN(n_2109));
   XOR2_X1 i_1910 (.A(n_2111), .B(n_2110), .Z(n_4156));
   NAND2_X1 i_1911 (.A1(inputB[28]), .A2(inputA[7]), .ZN(n_2110));
   OAI21_X1 i_1912 (.A(n_2112), .B1(n_2232), .B2(n_2114), .ZN(n_2111));
   NAND2_X1 i_1913 (.A1(n_2232), .A2(n_2114), .ZN(n_2112));
   INV_X1 i_1914 (.A(n_2115), .ZN(n_2114));
   NAND2_X1 i_1915 (.A1(inputB[26]), .A2(inputA[9]), .ZN(n_2115));
   XOR2_X1 i_1916 (.A(n_2117), .B(n_2116), .Z(n_4170));
   NAND2_X1 i_1917 (.A1(inputB[22]), .A2(inputA[13]), .ZN(n_2116));
   NAND2_X1 i_1918 (.A1(n_2119), .A2(n_2118), .ZN(n_2117));
   NAND3_X1 i_1919 (.A1(inputB[21]), .A2(inputA[14]), .A3(n_2123), .ZN(n_2118));
   INV_X1 i_1920 (.A(n_2122), .ZN(n_2119));
   AOI21_X1 i_1921 (.A(n_2123), .B1(inputB[21]), .B2(inputA[14]), .ZN(n_2122));
   AND2_X1 i_1922 (.A1(inputB[20]), .A2(inputA[15]), .ZN(n_2123));
   XOR2_X1 i_1923 (.A(n_2125), .B(n_2124), .Z(n_4177));
   NAND2_X1 i_1924 (.A1(inputB[19]), .A2(inputA[16]), .ZN(n_2124));
   NAND2_X1 i_1925 (.A1(n_2127), .A2(n_2126), .ZN(n_2125));
   NAND3_X1 i_1926 (.A1(inputB[17]), .A2(inputA[18]), .A3(n_2223), .ZN(n_2126));
   INV_X1 i_1927 (.A(n_2129), .ZN(n_2127));
   AOI21_X1 i_1928 (.A(n_2223), .B1(inputB[17]), .B2(inputA[18]), .ZN(n_2129));
   XOR2_X1 i_1929 (.A(n_2131), .B(n_2130), .Z(n_4191));
   NAND2_X1 i_1930 (.A1(inputB[13]), .A2(inputA[22]), .ZN(n_2130));
   NAND2_X1 i_1931 (.A1(n_2133), .A2(n_2132), .ZN(n_2131));
   NAND3_X1 i_1932 (.A1(inputB[12]), .A2(inputA[23]), .A3(n_2136), .ZN(n_2132));
   INV_X1 i_1933 (.A(n_2135), .ZN(n_2133));
   AOI21_X1 i_1934 (.A(n_2136), .B1(inputB[12]), .B2(inputA[23]), .ZN(n_2135));
   AND2_X1 i_1935 (.A1(inputB[11]), .A2(inputA[24]), .ZN(n_2136));
   XOR2_X1 i_1936 (.A(n_2138), .B(n_2137), .Z(n_4198));
   NAND2_X1 i_1938 (.A1(inputB[10]), .A2(inputA[25]), .ZN(n_2137));
   NAND2_X1 i_1939 (.A1(n_2140), .A2(n_2139), .ZN(n_2138));
   NAND4_X1 i_1940 (.A1(inputB[8]), .A2(inputA[26]), .A3(inputB[9]), .A4(
      inputA[27]), .ZN(n_2139));
   INV_X1 i_1942 (.A(n_2143), .ZN(n_2140));
   AOI22_X1 i_1943 (.A1(inputB[9]), .A2(inputA[26]), .B1(inputB[8]), .B2(
      inputA[27]), .ZN(n_2143));
   AOI21_X1 i_1944 (.A(n_2325), .B1(n_2324), .B2(n_2313), .ZN(n_4051));
   INV_X1 i_1946 (.A(n_2144), .ZN(n_4060));
   AOI21_X1 i_1947 (.A(n_4057), .B1(n_4056), .B2(n_2239), .ZN(n_2144));
   INV_X1 i_1948 (.A(n_2145), .ZN(n_4070));
   AOI21_X1 i_1950 (.A(n_4067), .B1(n_4066), .B2(n_2214), .ZN(n_2145));
   OAI21_X1 i_1951 (.A(n_2245), .B1(n_2252), .B2(n_2251), .ZN(n_3986));
   AOI22_X1 i_1952 (.A1(n_2446), .A2(n_2258), .B1(n_2256), .B2(n_2253), .ZN(
      n_4002));
   OAI21_X1 i_1954 (.A(n_2264), .B1(n_2268), .B2(n_2259), .ZN(n_4009));
   AOI21_X1 i_1955 (.A(n_2146), .B1(n_2456), .B2(n_2284), .ZN(n_4023));
   NOR2_X1 i_1956 (.A1(n_2279), .A2(n_2269), .ZN(n_2146));
   OAI21_X1 i_1958 (.A(n_2289), .B1(n_2299), .B2(n_2285), .ZN(n_4030));
   AOI22_X1 i_1959 (.A1(n_2466), .A2(n_2309), .B1(n_2304), .B2(n_2300), .ZN(
      n_4044));
   NAND2_X1 i_1960 (.A1(inputB[4]), .A2(inputA[31]), .ZN(n_384));
   INV_X1 i_1962 (.A(n_2150), .ZN(n_3978));
   AOI21_X1 i_1963 (.A(n_3975), .B1(n_3974), .B2(n_2154), .ZN(n_2150));
   INV_X1 i_1964 (.A(n_2155), .ZN(n_2154));
   AOI21_X1 i_1966 (.A(n_3803), .B1(n_3802), .B2(n_2474), .ZN(n_2155));
   XNOR2_X1 i_1967 (.A(n_4131), .B(n_2160), .ZN(n_4133));
   INV_X1 i_1968 (.A(n_2160), .ZN(n_2159));
   AOI21_X1 i_1970 (.A(n_3965), .B1(n_3964), .B2(n_2338), .ZN(n_2160));
   XNOR2_X1 i_1971 (.A(n_4126), .B(n_2165), .ZN(n_4128));
   INV_X1 i_1972 (.A(n_2165), .ZN(n_2161));
   AOI21_X1 i_1974 (.A(n_3955), .B1(n_3954), .B2(n_2335), .ZN(n_2165));
   XNOR2_X1 i_1975 (.A(n_4121), .B(n_2171), .ZN(n_4123));
   INV_X1 i_1976 (.A(n_2171), .ZN(n_2170));
   AOI21_X1 i_1978 (.A(n_3950), .B1(n_3949), .B2(n_2345), .ZN(n_2171));
   XNOR2_X1 i_1979 (.A(n_4116), .B(n_2175), .ZN(n_4118));
   INV_X1 i_1980 (.A(n_2175), .ZN(n_2174));
   AOI21_X1 i_1982 (.A(n_3940), .B1(n_3939), .B2(n_2362), .ZN(n_2175));
   XOR2_X1 i_1983 (.A(n_4111), .B(n_2180), .Z(n_4113));
   XOR2_X1 i_1984 (.A(n_4076), .B(n_2184), .Z(n_2180));
   XOR2_X1 i_1985 (.A(n_2186), .B(n_2185), .Z(n_2184));
   NAND2_X1 i_1986 (.A1(inputB[10]), .A2(inputA[24]), .ZN(n_2185));
   OAI21_X1 i_1987 (.A(n_2194), .B1(n_2460), .B2(n_2195), .ZN(n_2186));
   INV_X1 i_1988 (.A(n_2194), .ZN(n_2190));
   NAND2_X1 i_1989 (.A1(n_2460), .A2(n_2195), .ZN(n_2194));
   NAND2_X1 i_1990 (.A1(inputB[8]), .A2(inputA[26]), .ZN(n_2195));
   INV_X1 i_1991 (.A(n_2200), .ZN(n_3963));
   AOI21_X1 i_1992 (.A(n_3960), .B1(n_3959), .B2(n_2343), .ZN(n_2200));
   XNOR2_X1 i_1993 (.A(n_4106), .B(n_2205), .ZN(n_4108));
   INV_X1 i_1994 (.A(n_2205), .ZN(n_2204));
   AOI21_X1 i_1995 (.A(n_3930), .B1(n_3929), .B2(n_2358), .ZN(n_2205));
   XNOR2_X1 i_1996 (.A(n_4096), .B(n_2209), .ZN(n_4098));
   INV_X1 i_1997 (.A(n_2209), .ZN(n_2208));
   AOI21_X1 i_1998 (.A(n_3925), .B1(n_3924), .B2(n_2375), .ZN(n_2209));
   XNOR2_X1 i_1999 (.A(n_4101), .B(n_2211), .ZN(n_4103));
   INV_X1 i_2000 (.A(n_2211), .ZN(n_2210));
   AOI21_X1 i_2001 (.A(n_3910), .B1(n_3909), .B2(n_2363), .ZN(n_2211));
   INV_X1 i_2002 (.A(n_2212), .ZN(n_3948));
   AOI21_X1 i_2003 (.A(n_3945), .B1(n_3944), .B2(n_2355), .ZN(n_2212));
   XOR2_X1 i_2004 (.A(n_4091), .B(n_2213), .Z(n_4093));
   XOR2_X1 i_2005 (.A(n_4066), .B(n_2214), .Z(n_2213));
   AOI21_X1 i_2006 (.A(n_2391), .B1(n_2382), .B2(n_2376), .ZN(n_2214));
   XOR2_X1 i_2007 (.A(n_4081), .B(n_2215), .Z(n_4083));
   XOR2_X1 i_2008 (.A(n_2217), .B(n_2216), .Z(n_2215));
   NAND2_X1 i_2009 (.A1(inputB[19]), .A2(inputA[15]), .ZN(n_2216));
   NAND2_X1 i_2010 (.A1(n_2222), .A2(n_2218), .ZN(n_2217));
   INV_X1 i_2011 (.A(n_2219), .ZN(n_2218));
   AOI22_X1 i_2012 (.A1(inputB[18]), .A2(inputA[16]), .B1(inputB[17]), .B2(
      inputA[17]), .ZN(n_2219));
   NAND3_X1 i_2013 (.A1(inputB[17]), .A2(inputA[16]), .A3(n_2223), .ZN(n_2222));
   AND2_X1 i_2014 (.A1(inputB[18]), .A2(inputA[17]), .ZN(n_2223));
   XOR2_X1 i_2015 (.A(n_4086), .B(n_2224), .Z(n_4088));
   XOR2_X1 i_2016 (.A(n_2226), .B(n_2225), .Z(n_2224));
   NAND2_X1 i_2017 (.A1(inputB[28]), .A2(inputA[6]), .ZN(n_2225));
   NAND2_X1 i_2018 (.A1(n_2231), .A2(n_2229), .ZN(n_2226));
   INV_X1 i_2019 (.A(n_2230), .ZN(n_2229));
   AOI22_X1 i_2020 (.A1(inputB[27]), .A2(inputA[7]), .B1(inputB[26]), .B2(
      inputA[8]), .ZN(n_2230));
   NAND3_X1 i_2021 (.A1(inputB[26]), .A2(inputA[7]), .A3(n_2232), .ZN(n_2231));
   INV_X1 i_2022 (.A(n_2233), .ZN(n_2232));
   NAND2_X1 i_2023 (.A1(inputB[27]), .A2(inputA[8]), .ZN(n_2233));
   INV_X1 i_2024 (.A(n_2234), .ZN(n_3938));
   AOI21_X1 i_2025 (.A(n_3935), .B1(n_3934), .B2(n_2336), .ZN(n_2234));
   XNOR2_X1 i_2026 (.A(n_4071), .B(n_2236), .ZN(n_4073));
   INV_X1 i_2027 (.A(n_2236), .ZN(n_2235));
   AOI21_X1 i_2028 (.A(n_3890), .B1(n_3889), .B2(n_2412), .ZN(n_2236));
   INV_X1 i_2029 (.A(n_2237), .ZN(n_3918));
   AOI21_X1 i_2030 (.A(n_3915), .B1(n_3914), .B2(n_2346), .ZN(n_2237));
   INV_X1 i_2031 (.A(n_2238), .ZN(n_3923));
   AOI21_X1 i_2032 (.A(n_3920), .B1(n_3919), .B2(n_2369), .ZN(n_2238));
   XOR2_X1 i_2033 (.A(n_4056), .B(n_2239), .Z(n_4058));
   AOI21_X1 i_2034 (.A(n_2349), .B1(n_2524), .B2(n_2350), .ZN(n_2239));
   XOR2_X1 i_2035 (.A(n_4061), .B(n_2240), .Z(n_4063));
   OAI21_X1 i_2036 (.A(n_2372), .B1(n_2548), .B2(n_2371), .ZN(n_2240));
   INV_X1 i_2037 (.A(n_2243), .ZN(n_3908));
   AOI21_X1 i_2038 (.A(n_3905), .B1(n_3904), .B2(n_2397), .ZN(n_2243));
   XOR2_X1 i_2040 (.A(n_2252), .B(n_2244), .Z(n_3985));
   NAND2_X1 i_2041 (.A1(n_2250), .A2(n_2245), .ZN(n_2244));
   NAND3_X1 i_2042 (.A1(inputB[29]), .A2(inputA[4]), .A3(n_2246), .ZN(n_2245));
   INV_X1 i_2044 (.A(n_2247), .ZN(n_2246));
   NAND2_X1 i_2045 (.A1(inputB[30]), .A2(inputA[5]), .ZN(n_2247));
   INV_X1 i_2046 (.A(n_2251), .ZN(n_2250));
   AOI22_X1 i_2048 (.A1(inputB[30]), .A2(inputA[4]), .B1(inputB[29]), .B2(
      inputA[5]), .ZN(n_2251));
   AND2_X1 i_2049 (.A1(inputB[31]), .A2(inputA[3]), .ZN(n_2252));
   XNOR2_X1 i_2050 (.A(n_2254), .B(n_2253), .ZN(n_4001));
   NAND2_X1 i_2052 (.A1(inputB[25]), .A2(inputA[9]), .ZN(n_2253));
   AOI21_X1 i_2053 (.A(n_2257), .B1(n_2446), .B2(n_2258), .ZN(n_2254));
   INV_X1 i_2054 (.A(n_2257), .ZN(n_2256));
   NOR2_X1 i_2056 (.A1(n_2446), .A2(n_2258), .ZN(n_2257));
   NAND2_X1 i_2057 (.A1(inputB[23]), .A2(inputA[11]), .ZN(n_2258));
   XOR2_X1 i_2058 (.A(n_2260), .B(n_2259), .Z(n_4008));
   NAND2_X1 i_2060 (.A1(inputB[22]), .A2(inputA[12]), .ZN(n_2259));
   NAND2_X1 i_2061 (.A1(n_2265), .A2(n_2264), .ZN(n_2260));
   NAND3_X1 i_2062 (.A1(inputB[20]), .A2(inputA[14]), .A3(n_2373), .ZN(n_2264));
   INV_X1 i_2064 (.A(n_2268), .ZN(n_2265));
   AOI21_X1 i_2065 (.A(n_2373), .B1(inputB[20]), .B2(inputA[14]), .ZN(n_2268));
   XOR2_X1 i_2066 (.A(n_2274), .B(n_2269), .Z(n_4022));
   AND2_X1 i_2068 (.A1(inputB[16]), .A2(inputA[18]), .ZN(n_2269));
   AOI21_X1 i_2069 (.A(n_2279), .B1(n_2456), .B2(n_2284), .ZN(n_2274));
   NOR2_X1 i_2070 (.A1(n_2456), .A2(n_2284), .ZN(n_2279));
   NAND2_X1 i_2072 (.A1(inputB[14]), .A2(inputA[20]), .ZN(n_2284));
   XOR2_X1 i_2073 (.A(n_2288), .B(n_2285), .Z(n_4029));
   NAND2_X1 i_2074 (.A1(inputB[13]), .A2(inputA[21]), .ZN(n_2285));
   NAND2_X1 i_2076 (.A1(n_2294), .A2(n_2289), .ZN(n_2288));
   NAND3_X1 i_2077 (.A1(inputB[11]), .A2(inputA[23]), .A3(n_2351), .ZN(n_2289));
   INV_X1 i_2078 (.A(n_2299), .ZN(n_2294));
   AOI21_X1 i_2080 (.A(n_2351), .B1(inputB[11]), .B2(inputA[23]), .ZN(n_2299));
   XNOR2_X1 i_2081 (.A(n_2303), .B(n_2300), .ZN(n_4043));
   NAND2_X1 i_2082 (.A1(inputB[7]), .A2(inputA[27]), .ZN(n_2300));
   AOI21_X1 i_2084 (.A(n_2305), .B1(n_2466), .B2(n_2309), .ZN(n_2303));
   INV_X1 i_2085 (.A(n_2305), .ZN(n_2304));
   NOR2_X1 i_2086 (.A1(n_2466), .A2(n_2309), .ZN(n_2305));
   NAND2_X1 i_2087 (.A1(inputB[5]), .A2(inputA[29]), .ZN(n_2309));
   XOR2_X1 i_2088 (.A(n_2319), .B(n_2314), .Z(n_4050));
   INV_X1 i_2089 (.A(n_2314), .ZN(n_2313));
   AOI21_X1 i_2090 (.A(n_2367), .B1(n_2487), .B2(n_2365), .ZN(n_2314));
   NOR2_X1 i_2091 (.A1(n_2325), .A2(n_2323), .ZN(n_2319));
   INV_X1 i_2092 (.A(n_2324), .ZN(n_2323));
   OAI211_X1 i_2093 (.A(inputB[4]), .B(inputA[30]), .C1(n_5756), .C2(n_5753), 
      .ZN(n_2324));
   AOI211_X1 i_2094 (.A(n_5756), .B(n_5753), .C1(inputB[4]), .C2(inputA[30]), 
      .ZN(n_2325));
   INV_X1 i_2095 (.A(n_2326), .ZN(n_3898));
   AOI21_X1 i_2096 (.A(n_3895), .B1(n_3894), .B2(n_2359), .ZN(n_2326));
   INV_X1 i_2097 (.A(n_2327), .ZN(n_3903));
   AOI21_X1 i_2098 (.A(n_3900), .B1(n_3899), .B2(n_2417), .ZN(n_2327));
   OAI21_X1 i_2099 (.A(n_2427), .B1(n_2585), .B2(n_2432), .ZN(n_3828));
   NOR2_X1 i_2100 (.A1(n_2437), .A2(n_2328), .ZN(n_3835));
   NOR2_X1 i_2101 (.A1(n_2590), .A2(n_2442), .ZN(n_2328));
   OAI21_X1 i_2102 (.A(n_2450), .B1(n_2603), .B2(n_2452), .ZN(n_3849));
   NOR2_X1 i_2103 (.A1(n_2454), .A2(n_2329), .ZN(n_3856));
   NOR2_X1 i_2104 (.A1(n_2607), .A2(n_2455), .ZN(n_2329));
   NOR2_X1 i_2105 (.A1(n_2458), .A2(n_2330), .ZN(n_3870));
   NOR2_X1 i_2106 (.A1(n_2618), .A2(n_2459), .ZN(n_2330));
   OAI22_X1 i_2107 (.A1(n_2481), .A2(n_2466), .B1(n_2625), .B2(n_2464), .ZN(
      n_3877));
   INV_X1 i_2108 (.A(n_2331), .ZN(n_3811));
   AOI21_X1 i_2109 (.A(n_3808), .B1(n_3807), .B2(n_2472), .ZN(n_2331));
   XOR2_X1 i_2110 (.A(n_3969), .B(n_2334), .Z(n_3971));
   XOR2_X1 i_2111 (.A(n_3954), .B(n_2335), .Z(n_2334));
   XNOR2_X1 i_2112 (.A(n_3934), .B(n_2337), .ZN(n_2335));
   INV_X1 i_2113 (.A(n_2337), .ZN(n_2336));
   AOI21_X1 i_2114 (.A(n_3753), .B1(n_3752), .B2(n_2527), .ZN(n_2337));
   XNOR2_X1 i_2115 (.A(n_3964), .B(n_2341), .ZN(n_3966));
   INV_X1 i_2116 (.A(n_2341), .ZN(n_2338));
   AOI21_X1 i_2117 (.A(n_3793), .B1(n_3792), .B2(n_2475), .ZN(n_2341));
   INV_X1 i_2118 (.A(n_2342), .ZN(n_3801));
   AOI21_X1 i_2119 (.A(n_3798), .B1(n_3797), .B2(n_2477), .ZN(n_2342));
   XNOR2_X1 i_2120 (.A(n_3959), .B(n_2344), .ZN(n_3961));
   INV_X1 i_2121 (.A(n_2344), .ZN(n_2343));
   AOI21_X1 i_2122 (.A(n_3778), .B1(n_3777), .B2(n_2497), .ZN(n_2344));
   XOR2_X1 i_2123 (.A(n_3949), .B(n_2345), .Z(n_3951));
   XOR2_X1 i_2124 (.A(n_3914), .B(n_2346), .Z(n_2345));
   XNOR2_X1 i_2125 (.A(n_2523), .B(n_2347), .ZN(n_2346));
   NAND2_X1 i_2126 (.A1(n_2350), .A2(n_2348), .ZN(n_2347));
   INV_X1 i_2127 (.A(n_2349), .ZN(n_2348));
   AOI22_X1 i_2128 (.A1(inputB[11]), .A2(inputA[22]), .B1(inputB[12]), .B2(
      inputA[21]), .ZN(n_2349));
   NAND3_X1 i_2129 (.A1(inputB[11]), .A2(inputA[21]), .A3(n_2351), .ZN(n_2350));
   AND2_X1 i_2130 (.A1(inputB[12]), .A2(inputA[22]), .ZN(n_2351));
   INV_X1 i_2131 (.A(n_2352), .ZN(n_3791));
   AOI21_X1 i_2132 (.A(n_3788), .B1(n_3787), .B2(n_2489), .ZN(n_2352));
   XNOR2_X1 i_2133 (.A(n_3944), .B(n_2356), .ZN(n_3946));
   INV_X1 i_2134 (.A(n_2356), .ZN(n_2355));
   AOI21_X1 i_2135 (.A(n_3763), .B1(n_3762), .B2(n_2492), .ZN(n_2356));
   INV_X1 i_2136 (.A(n_2357), .ZN(n_3786));
   AOI21_X1 i_2137 (.A(n_3783), .B1(n_3782), .B2(n_2478), .ZN(n_2357));
   XOR2_X1 i_2138 (.A(n_3929), .B(n_2358), .Z(n_3931));
   XOR2_X1 i_2139 (.A(n_3894), .B(n_2359), .Z(n_2358));
   AOI21_X1 i_2140 (.A(n_2598), .B1(n_2599), .B2(n_2595), .ZN(n_2359));
   XOR2_X1 i_2142 (.A(n_3939), .B(n_2362), .Z(n_3941));
   XOR2_X1 i_2143 (.A(n_3909), .B(n_2363), .Z(n_2362));
   XOR2_X1 i_2144 (.A(n_2487), .B(n_2364), .Z(n_2363));
   NAND2_X1 i_2146 (.A1(n_2366), .A2(n_2365), .ZN(n_2364));
   OAI211_X1 i_2147 (.A(inputB[3]), .B(inputA[30]), .C1(n_5755), .C2(n_5753), 
      .ZN(n_2365));
   INV_X1 i_2148 (.A(n_2367), .ZN(n_2366));
   AOI211_X1 i_2150 (.A(n_5755), .B(n_5753), .C1(inputB[3]), .C2(inputA[30]), 
      .ZN(n_2367));
   INV_X1 i_2151 (.A(n_2368), .ZN(n_3776));
   AOI21_X1 i_2152 (.A(n_3773), .B1(n_3772), .B2(n_2500), .ZN(n_2368));
   XOR2_X1 i_2154 (.A(n_3919), .B(n_2369), .Z(n_3921));
   XOR2_X1 i_2155 (.A(n_2547), .B(n_2370), .Z(n_2369));
   AOI21_X1 i_2156 (.A(n_2371), .B1(n_2594), .B2(n_2373), .ZN(n_2370));
   AOI22_X1 i_2158 (.A1(inputB[20]), .A2(inputA[13]), .B1(inputB[21]), .B2(
      inputA[12]), .ZN(n_2371));
   NAND2_X1 i_2159 (.A1(n_2594), .A2(n_2373), .ZN(n_2372));
   AND2_X1 i_2160 (.A1(inputB[21]), .A2(inputA[13]), .ZN(n_2373));
   XOR2_X1 i_2162 (.A(n_3924), .B(n_2375), .Z(n_3926));
   XNOR2_X1 i_2163 (.A(n_2378), .B(n_2377), .ZN(n_2375));
   INV_X1 i_2164 (.A(n_2377), .ZN(n_2376));
   NAND2_X1 i_2166 (.A1(inputB[31]), .A2(inputA[2]), .ZN(n_2377));
   NAND2_X1 i_2167 (.A1(n_2387), .A2(n_2382), .ZN(n_2378));
   NAND4_X1 i_2168 (.A1(inputB[29]), .A2(inputA[3]), .A3(inputB[30]), .A4(
      inputA[4]), .ZN(n_2382));
   INV_X1 i_2170 (.A(n_2391), .ZN(n_2387));
   AOI22_X1 i_2171 (.A1(inputB[29]), .A2(inputA[4]), .B1(inputB[30]), .B2(
      inputA[3]), .ZN(n_2391));
   INV_X1 i_2172 (.A(n_2392), .ZN(n_3771));
   AOI21_X1 i_2174 (.A(n_3768), .B1(n_3767), .B2(n_2506), .ZN(n_2392));
   XNOR2_X1 i_2175 (.A(n_3904), .B(n_2402), .ZN(n_3906));
   INV_X1 i_2176 (.A(n_2402), .ZN(n_2397));
   AOI21_X1 i_2178 (.A(n_3728), .B1(n_3727), .B2(n_2493), .ZN(n_2402));
   INV_X1 i_2179 (.A(n_2406), .ZN(n_3746));
   AOI21_X1 i_2180 (.A(n_3743), .B1(n_3742), .B2(n_2479), .ZN(n_2406));
   INV_X1 i_2182 (.A(n_2407), .ZN(n_3751));
   AOI21_X1 i_2183 (.A(n_3748), .B1(n_3747), .B2(n_2509), .ZN(n_2407));
   INV_X1 i_2184 (.A(n_2408), .ZN(n_3761));
   AOI21_X1 i_2186 (.A(n_3758), .B1(n_3757), .B2(n_2498), .ZN(n_2408));
   XOR2_X1 i_2187 (.A(n_3889), .B(n_2412), .Z(n_3891));
   OAI21_X1 i_2188 (.A(n_2617), .B1(n_2616), .B2(n_2612), .ZN(n_2412));
   XOR2_X1 i_2190 (.A(n_3899), .B(n_2417), .Z(n_3901));
   OAI21_X1 i_2191 (.A(n_2583), .B1(n_2582), .B2(n_2577), .ZN(n_2417));
   INV_X1 i_2192 (.A(n_2422), .ZN(n_3741));
   AOI21_X1 i_2193 (.A(n_3738), .B1(n_3737), .B2(n_2501), .ZN(n_2422));
   XNOR2_X1 i_2194 (.A(n_2584), .B(n_2426), .ZN(n_3827));
   NAND2_X1 i_2195 (.A1(n_2428), .A2(n_2427), .ZN(n_2426));
   NAND4_X1 i_2196 (.A1(inputB[26]), .A2(inputA[7]), .A3(inputB[27]), .A4(
      inputA[6]), .ZN(n_2427));
   INV_X1 i_2197 (.A(n_2432), .ZN(n_2428));
   AOI22_X1 i_2198 (.A1(inputB[26]), .A2(inputA[7]), .B1(inputB[27]), .B2(
      inputA[6]), .ZN(n_2432));
   XOR2_X1 i_2199 (.A(n_2590), .B(n_2436), .Z(n_3834));
   NOR2_X1 i_2200 (.A1(n_2442), .A2(n_2437), .ZN(n_2436));
   AOI22_X1 i_2201 (.A1(inputB[23]), .A2(inputA[10]), .B1(inputB[24]), .B2(
      inputA[9]), .ZN(n_2437));
   NOR2_X1 i_2202 (.A1(n_2528), .A2(n_2446), .ZN(n_2442));
   NAND2_X1 i_2203 (.A1(inputB[24]), .A2(inputA[10]), .ZN(n_2446));
   XNOR2_X1 i_2204 (.A(n_2602), .B(n_2447), .ZN(n_3848));
   NAND2_X1 i_2205 (.A1(n_2451), .A2(n_2450), .ZN(n_2447));
   NAND3_X1 i_2206 (.A1(inputB[18]), .A2(inputA[16]), .A3(n_2610), .ZN(n_2450));
   INV_X1 i_2207 (.A(n_2452), .ZN(n_2451));
   AOI22_X1 i_2208 (.A1(inputB[17]), .A2(inputA[16]), .B1(inputB[18]), .B2(
      inputA[15]), .ZN(n_2452));
   XOR2_X1 i_2209 (.A(n_2607), .B(n_2453), .Z(n_3855));
   NOR2_X1 i_2210 (.A1(n_2455), .A2(n_2454), .ZN(n_2453));
   AOI22_X1 i_2211 (.A1(inputB[14]), .A2(inputA[19]), .B1(inputB[15]), .B2(
      inputA[18]), .ZN(n_2454));
   NOR2_X1 i_2212 (.A1(n_2513), .A2(n_2456), .ZN(n_2455));
   NAND2_X1 i_2213 (.A1(inputB[15]), .A2(inputA[19]), .ZN(n_2456));
   XOR2_X1 i_2214 (.A(n_2618), .B(n_2457), .Z(n_3869));
   NOR2_X1 i_2215 (.A1(n_2459), .A2(n_2458), .ZN(n_2457));
   AOI22_X1 i_2216 (.A1(inputB[8]), .A2(inputA[25]), .B1(inputB[9]), .B2(
      inputA[24]), .ZN(n_2458));
   NOR2_X1 i_2217 (.A1(n_2619), .A2(n_2460), .ZN(n_2459));
   NAND2_X1 i_2218 (.A1(inputB[9]), .A2(inputA[25]), .ZN(n_2460));
   XOR2_X1 i_2219 (.A(n_2624), .B(n_2461), .Z(n_3876));
   AOI21_X1 i_2220 (.A(n_2464), .B1(n_2480), .B2(n_2465), .ZN(n_2461));
   AOI22_X1 i_2221 (.A1(inputB[5]), .A2(inputA[28]), .B1(inputB[6]), .B2(
      inputA[27]), .ZN(n_2464));
   INV_X1 i_2222 (.A(n_2466), .ZN(n_2465));
   NAND2_X1 i_2223 (.A1(inputB[6]), .A2(inputA[28]), .ZN(n_2466));
   AND2_X1 i_2224 (.A1(n_2638), .A2(n_2631), .ZN(n_3717));
   INV_X1 i_2225 (.A(n_2467), .ZN(n_3726));
   AOI21_X1 i_2226 (.A(n_3723), .B1(n_3722), .B2(n_2567), .ZN(n_2467));
   INV_X1 i_2227 (.A(n_2468), .ZN(n_3736));
   AOI21_X1 i_2228 (.A(n_3733), .B1(n_3732), .B2(n_2568), .ZN(n_2468));
   OAI21_X1 i_2229 (.A(n_2589), .B1(n_2592), .B2(n_2586), .ZN(n_3661));
   OAI21_X1 i_2230 (.A(n_2543), .B1(n_2539), .B2(n_2528), .ZN(n_3668));
   OAI21_X1 i_2231 (.A(n_2606), .B1(n_2611), .B2(n_2609), .ZN(n_3682));
   OAI21_X1 i_2232 (.A(n_2522), .B1(n_2518), .B2(n_2513), .ZN(n_3689));
   OAI21_X1 i_2233 (.A(n_2623), .B1(n_2627), .B2(n_2619), .ZN(n_3703));
   OAI21_X1 i_2234 (.A(n_2471), .B1(n_2819), .B2(n_2487), .ZN(n_3710));
   NAND2_X1 i_2235 (.A1(n_2485), .A2(n_2480), .ZN(n_2471));
   XNOR2_X1 i_2236 (.A(n_3807), .B(n_2473), .ZN(n_3809));
   INV_X1 i_2237 (.A(n_2473), .ZN(n_2472));
   AOI21_X1 i_2238 (.A(n_3636), .B1(n_3635), .B2(n_2649), .ZN(n_2473));
   XOR2_X1 i_2239 (.A(n_3802), .B(n_2474), .Z(n_3804));
   XNOR2_X1 i_2240 (.A(n_3792), .B(n_2476), .ZN(n_2474));
   INV_X1 i_2241 (.A(n_2476), .ZN(n_2475));
   AOI21_X1 i_2242 (.A(n_3616), .B1(n_3615), .B2(n_2699), .ZN(n_2476));
   XOR2_X1 i_2243 (.A(n_3797), .B(n_2477), .Z(n_3799));
   XOR2_X1 i_2244 (.A(n_3782), .B(n_2478), .Z(n_2477));
   XOR2_X1 i_2245 (.A(n_3742), .B(n_2479), .Z(n_2478));
   XOR2_X1 i_2247 (.A(n_2482), .B(n_2481), .Z(n_2479));
   INV_X1 i_2248 (.A(n_2481), .ZN(n_2480));
   NAND2_X1 i_2249 (.A1(inputB[5]), .A2(inputA[27]), .ZN(n_2481));
   OAI21_X1 i_2251 (.A(n_2485), .B1(n_2819), .B2(n_2487), .ZN(n_2482));
   OAI21_X1 i_2252 (.A(n_2486), .B1(n_5756), .B2(n_5750), .ZN(n_2485));
   NAND2_X1 i_2253 (.A1(inputB[4]), .A2(inputA[28]), .ZN(n_2486));
   NAND2_X1 i_2255 (.A1(inputB[4]), .A2(inputA[29]), .ZN(n_2487));
   INV_X1 i_2256 (.A(n_2488), .ZN(n_3634));
   AOI21_X1 i_2257 (.A(n_3631), .B1(n_3630), .B2(n_2658), .ZN(n_2488));
   XOR2_X1 i_2259 (.A(n_3787), .B(n_2489), .Z(n_3789));
   XOR2_X1 i_2260 (.A(n_3762), .B(n_2492), .Z(n_2489));
   XOR2_X1 i_2261 (.A(n_3727), .B(n_2493), .Z(n_2492));
   NAND2_X1 i_2263 (.A1(n_2765), .A2(n_2494), .ZN(n_2493));
   NAND2_X1 i_2264 (.A1(n_2763), .A2(n_2761), .ZN(n_2494));
   INV_X1 i_2265 (.A(n_2495), .ZN(n_3629));
   AOI21_X1 i_2267 (.A(n_3626), .B1(n_3625), .B2(n_2650), .ZN(n_2495));
   INV_X1 i_2268 (.A(n_2496), .ZN(n_3624));
   AOI21_X1 i_2269 (.A(n_3621), .B1(n_3620), .B2(n_2669), .ZN(n_2496));
   XOR2_X1 i_2271 (.A(n_3777), .B(n_2497), .Z(n_3779));
   XOR2_X1 i_2272 (.A(n_3757), .B(n_2498), .Z(n_2497));
   OAI21_X1 i_2273 (.A(n_3649), .B1(n_2749), .B2(n_2499), .ZN(n_2498));
   NAND2_X1 i_2275 (.A1(n_2749), .A2(n_2499), .ZN(n_3649));
   AND2_X1 i_2276 (.A1(inputB[31]), .A2(inputA[1]), .ZN(n_2499));
   XOR2_X1 i_2277 (.A(n_3772), .B(n_2500), .Z(n_3774));
   XNOR2_X1 i_2279 (.A(n_3737), .B(n_2502), .ZN(n_2500));
   INV_X1 i_2280 (.A(n_2502), .ZN(n_2501));
   AOI21_X1 i_2281 (.A(n_3556), .B1(n_3555), .B2(n_2674), .ZN(n_2502));
   INV_X1 i_2283 (.A(n_2503), .ZN(n_3614));
   AOI21_X1 i_2284 (.A(n_3611), .B1(n_3610), .B2(n_2675), .ZN(n_2503));
   XNOR2_X1 i_2285 (.A(n_3767), .B(n_2507), .ZN(n_3769));
   INV_X1 i_2287 (.A(n_2507), .ZN(n_2506));
   AOI21_X1 i_2288 (.A(n_3581), .B1(n_3580), .B2(n_2726), .ZN(n_2507));
   INV_X1 i_2289 (.A(n_2508), .ZN(n_3609));
   AOI21_X1 i_2291 (.A(n_3606), .B1(n_3605), .B2(n_2704), .ZN(n_2508));
   XOR2_X1 i_2292 (.A(n_3747), .B(n_2509), .Z(n_3749));
   XOR2_X1 i_2293 (.A(n_2514), .B(n_2513), .Z(n_2509));
   NAND2_X1 i_2295 (.A1(inputB[14]), .A2(inputA[18]), .ZN(n_2513));
   NAND2_X1 i_2296 (.A1(n_2522), .A2(n_2517), .ZN(n_2514));
   INV_X1 i_2297 (.A(n_2518), .ZN(n_2517));
   AOI22_X1 i_2299 (.A1(inputB[12]), .A2(inputA[20]), .B1(inputB[13]), .B2(
      inputA[19]), .ZN(n_2518));
   NAND2_X1 i_2300 (.A1(n_2779), .A2(n_2523), .ZN(n_2522));
   INV_X1 i_2301 (.A(n_2524), .ZN(n_2523));
   NAND2_X1 i_2302 (.A1(inputB[13]), .A2(inputA[20]), .ZN(n_2524));
   XOR2_X1 i_2303 (.A(n_3752), .B(n_2527), .Z(n_3754));
   XOR2_X1 i_2304 (.A(n_2533), .B(n_2528), .Z(n_2527));
   NAND2_X1 i_2305 (.A1(inputB[23]), .A2(inputA[9]), .ZN(n_2528));
   NAND2_X1 i_2306 (.A1(n_2543), .A2(n_2538), .ZN(n_2533));
   INV_X1 i_2307 (.A(n_2539), .ZN(n_2538));
   AOI22_X1 i_2308 (.A1(inputB[21]), .A2(inputA[11]), .B1(inputB[22]), .B2(
      inputA[10]), .ZN(n_2539));
   NAND2_X1 i_2309 (.A1(n_2766), .A2(n_2547), .ZN(n_2543));
   INV_X1 i_2310 (.A(n_2548), .ZN(n_2547));
   NAND2_X1 i_2311 (.A1(inputB[22]), .A2(inputA[11]), .ZN(n_2548));
   INV_X1 i_2312 (.A(n_2553), .ZN(n_3599));
   AOI21_X1 i_2313 (.A(n_3596), .B1(n_3595), .B2(n_2673), .ZN(n_2553));
   INV_X1 i_2314 (.A(n_2557), .ZN(n_3604));
   AOI21_X1 i_2315 (.A(n_3601), .B1(n_3600), .B2(n_2714), .ZN(n_2557));
   INV_X1 i_2316 (.A(n_2558), .ZN(n_3594));
   AOI21_X1 i_2317 (.A(n_3591), .B1(n_3590), .B2(n_2733), .ZN(n_2558));
   INV_X1 i_2318 (.A(n_2559), .ZN(n_3579));
   AOI21_X1 i_2319 (.A(n_3576), .B1(n_3575), .B2(n_2719), .ZN(n_2559));
   INV_X1 i_2320 (.A(n_2563), .ZN(n_3589));
   AOI21_X1 i_2321 (.A(n_3586), .B1(n_3585), .B2(n_2679), .ZN(n_2563));
   XOR2_X1 i_2322 (.A(n_3722), .B(n_2567), .Z(n_3724));
   AOI22_X1 i_2323 (.A1(n_2872), .A2(n_2780), .B1(n_2778), .B2(n_2774), .ZN(
      n_2567));
   XOR2_X1 i_2324 (.A(n_3732), .B(n_2568), .Z(n_3734));
   AOI21_X1 i_2325 (.A(n_2752), .B1(n_2748), .B2(n_2745), .ZN(n_2568));
   INV_X1 i_2326 (.A(n_2573), .ZN(n_3574));
   AOI21_X1 i_2327 (.A(n_3571), .B1(n_3570), .B2(n_2738), .ZN(n_2573));
   XOR2_X1 i_2328 (.A(n_2578), .B(n_2577), .Z(n_3653));
   NAND2_X1 i_2329 (.A1(inputB[29]), .A2(inputA[3]), .ZN(n_2577));
   NAND2_X1 i_2330 (.A1(n_2583), .A2(n_2581), .ZN(n_2578));
   INV_X1 i_2331 (.A(n_2582), .ZN(n_2581));
   AOI22_X1 i_2332 (.A1(inputB[27]), .A2(inputA[5]), .B1(inputB[28]), .B2(
      inputA[4]), .ZN(n_2582));
   NAND2_X1 i_2333 (.A1(n_2760), .A2(n_2584), .ZN(n_2583));
   INV_X1 i_2334 (.A(n_2585), .ZN(n_2584));
   NAND2_X1 i_2335 (.A1(inputB[28]), .A2(inputA[5]), .ZN(n_2585));
   XOR2_X1 i_2336 (.A(n_2588), .B(n_2586), .Z(n_3660));
   NAND2_X1 i_2337 (.A1(inputB[26]), .A2(inputA[6]), .ZN(n_2586));
   NAND2_X1 i_2338 (.A1(n_2591), .A2(n_2589), .ZN(n_2588));
   NAND3_X1 i_2339 (.A1(inputB[24]), .A2(inputA[7]), .A3(n_2590), .ZN(n_2589));
   AND2_X1 i_2340 (.A1(inputB[25]), .A2(inputA[8]), .ZN(n_2590));
   INV_X1 i_2341 (.A(n_2592), .ZN(n_2591));
   AOI22_X1 i_2342 (.A1(inputB[24]), .A2(inputA[8]), .B1(inputB[25]), .B2(
      inputA[7]), .ZN(n_2592));
   XNOR2_X1 i_2343 (.A(n_2596), .B(n_2594), .ZN(n_3674));
   INV_X1 i_2344 (.A(n_2595), .ZN(n_2594));
   NAND2_X1 i_2345 (.A1(inputB[20]), .A2(inputA[12]), .ZN(n_2595));
   NAND2_X1 i_2346 (.A1(n_2599), .A2(n_2597), .ZN(n_2596));
   INV_X1 i_2347 (.A(n_2598), .ZN(n_2597));
   AOI22_X1 i_2348 (.A1(inputB[18]), .A2(inputA[14]), .B1(inputB[19]), .B2(
      inputA[13]), .ZN(n_2598));
   NAND2_X1 i_2349 (.A1(n_2773), .A2(n_2602), .ZN(n_2599));
   INV_X1 i_2350 (.A(n_2603), .ZN(n_2602));
   NAND2_X1 i_2351 (.A1(inputB[19]), .A2(inputA[14]), .ZN(n_2603));
   XOR2_X1 i_2352 (.A(n_2610), .B(n_2604), .Z(n_3681));
   NOR2_X1 i_2353 (.A1(n_2609), .A2(n_2605), .ZN(n_2604));
   INV_X1 i_2354 (.A(n_2606), .ZN(n_2605));
   NAND3_X1 i_2355 (.A1(inputB[15]), .A2(inputA[16]), .A3(n_2607), .ZN(n_2606));
   AND2_X1 i_2356 (.A1(inputB[16]), .A2(inputA[17]), .ZN(n_2607));
   AOI22_X1 i_2357 (.A1(inputB[15]), .A2(inputA[17]), .B1(inputB[16]), .B2(
      inputA[16]), .ZN(n_2609));
   INV_X1 i_2358 (.A(n_2611), .ZN(n_2610));
   NAND2_X1 i_2359 (.A1(inputB[17]), .A2(inputA[15]), .ZN(n_2611));
   XOR2_X1 i_2360 (.A(n_2613), .B(n_2612), .Z(n_3695));
   NAND2_X1 i_2361 (.A1(inputB[11]), .A2(inputA[21]), .ZN(n_2612));
   NAND2_X1 i_2362 (.A1(n_2617), .A2(n_2615), .ZN(n_2613));
   INV_X1 i_2364 (.A(n_2616), .ZN(n_2615));
   AOI22_X1 i_2365 (.A1(inputB[9]), .A2(inputA[23]), .B1(inputB[10]), .B2(
      inputA[22]), .ZN(n_2616));
   NAND2_X1 i_2366 (.A1(n_2800), .A2(n_2618), .ZN(n_2617));
   AND2_X1 i_2368 (.A1(inputB[10]), .A2(inputA[23]), .ZN(n_2618));
   XOR2_X1 i_2369 (.A(n_2620), .B(n_2619), .Z(n_3702));
   NAND2_X1 i_2370 (.A1(inputB[8]), .A2(inputA[24]), .ZN(n_2619));
   NAND2_X1 i_2372 (.A1(n_2626), .A2(n_2623), .ZN(n_2620));
   NAND3_X1 i_2373 (.A1(inputB[6]), .A2(inputA[25]), .A3(n_2624), .ZN(n_2623));
   INV_X1 i_2374 (.A(n_2625), .ZN(n_2624));
   NAND2_X1 i_2376 (.A1(inputB[7]), .A2(inputA[26]), .ZN(n_2625));
   INV_X1 i_2377 (.A(n_2627), .ZN(n_2626));
   AOI22_X1 i_2378 (.A1(inputB[6]), .A2(inputA[26]), .B1(inputB[7]), .B2(
      inputA[25]), .ZN(n_2627));
   INV_X1 i_2380 (.A(n_2628), .ZN(n_3716));
   AOI21_X1 i_2381 (.A(n_2632), .B1(n_2638), .B2(n_2630), .ZN(n_2628));
   INV_X1 i_2382 (.A(n_2631), .ZN(n_2630));
   NAND2_X1 i_2384 (.A1(n_2637), .A2(n_2633), .ZN(n_2631));
   AOI21_X1 i_2385 (.A(n_2633), .B1(n_2638), .B2(n_2637), .ZN(n_2632));
   NAND2_X1 i_2386 (.A1(n_2813), .A2(n_2636), .ZN(n_2633));
   NAND2_X1 i_2388 (.A1(n_2814), .A2(n_2804), .ZN(n_2636));
   OAI211_X1 i_2389 (.A(inputB[2]), .B(inputA[30]), .C1(n_5754), .C2(n_5753), 
      .ZN(n_2637));
   OAI211_X1 i_2390 (.A(inputB[1]), .B(inputA[31]), .C1(n_5755), .C2(n_5751), 
      .ZN(n_2638));
   INV_X1 i_2392 (.A(n_2639), .ZN(n_3550));
   AOI21_X1 i_2393 (.A(n_2830), .B1(n_2833), .B2(n_2824), .ZN(n_2639));
   INV_X1 i_2394 (.A(n_2640), .ZN(n_3564));
   AOI21_X1 i_2396 (.A(n_3561), .B1(n_3560), .B2(n_2742), .ZN(n_2640));
   INV_X1 i_2397 (.A(n_2643), .ZN(n_3569));
   AOI21_X1 i_2398 (.A(n_3566), .B1(n_3565), .B2(n_2744), .ZN(n_2643));
   OAI21_X1 i_2400 (.A(n_2755), .B1(n_2759), .B2(n_2753), .ZN(n_3487));
   OAI21_X1 i_2401 (.A(n_2695), .B1(n_2694), .B2(n_2684), .ZN(n_3494));
   OAI21_X1 i_2402 (.A(n_2770), .B1(n_2772), .B2(n_2768), .ZN(n_3508));
   OAI21_X1 i_2404 (.A(n_2732), .B1(n_2731), .B2(n_2727), .ZN(n_3515));
   OAI21_X1 i_2405 (.A(n_2794), .B1(n_2799), .B2(n_2784), .ZN(n_3529));
   OAI21_X1 i_2406 (.A(n_2725), .B1(n_2724), .B2(n_2720), .ZN(n_3536));
   XOR2_X1 i_2408 (.A(n_3640), .B(n_2644), .Z(n_3642));
   XOR2_X1 i_2409 (.A(n_3635), .B(n_2649), .Z(n_2644));
   XNOR2_X1 i_2410 (.A(n_3625), .B(n_2654), .ZN(n_2649));
   INV_X1 i_2412 (.A(n_2654), .ZN(n_2650));
   AOI21_X1 i_2413 (.A(n_3450), .B1(n_3449), .B2(n_2857), .ZN(n_2654));
   INV_X1 i_2414 (.A(n_2655), .ZN(n_3473));
   AOI21_X1 i_2416 (.A(n_3470), .B1(n_3469), .B2(n_2839), .ZN(n_2655));
   XNOR2_X1 i_2417 (.A(n_3630), .B(n_2659), .ZN(n_3632));
   INV_X1 i_2418 (.A(n_2659), .ZN(n_2658));
   AOI21_X1 i_2419 (.A(n_3455), .B1(n_3454), .B2(n_2860), .ZN(n_2659));
   INV_X1 i_2420 (.A(n_2660), .ZN(n_3468));
   AOI21_X1 i_2421 (.A(n_3465), .B1(n_3464), .B2(n_2843), .ZN(n_2660));
   INV_X1 i_2422 (.A(n_2664), .ZN(n_3463));
   AOI21_X1 i_2423 (.A(n_3460), .B1(n_3459), .B2(n_2853), .ZN(n_2664));
   XOR2_X1 i_2424 (.A(n_3620), .B(n_2669), .Z(n_3622));
   XOR2_X1 i_2425 (.A(n_3595), .B(n_2673), .Z(n_2669));
   XOR2_X1 i_2426 (.A(n_3555), .B(n_2674), .Z(n_2673));
   OAI21_X1 i_2427 (.A(n_2870), .B1(n_2874), .B2(n_2867), .ZN(n_2674));
   XOR2_X1 i_2428 (.A(n_3610), .B(n_2675), .Z(n_3612));
   XOR2_X1 i_2429 (.A(n_3585), .B(n_2679), .Z(n_2675));
   XOR2_X1 i_2430 (.A(n_2689), .B(n_2684), .Z(n_2679));
   NAND2_X1 i_2431 (.A1(inputB[25]), .A2(inputA[6]), .ZN(n_2684));
   NAND2_X1 i_2432 (.A1(n_2695), .A2(n_2693), .ZN(n_2689));
   INV_X1 i_2433 (.A(n_2694), .ZN(n_2693));
   AOI22_X1 i_2434 (.A1(inputB[23]), .A2(inputA[8]), .B1(inputB[24]), .B2(
      inputA[7]), .ZN(n_2694));
   NAND3_X1 i_2435 (.A1(inputB[24]), .A2(inputA[8]), .A3(n_2962), .ZN(n_2695));
   XNOR2_X1 i_2436 (.A(n_3615), .B(n_2703), .ZN(n_3617));
   INV_X1 i_2437 (.A(n_2703), .ZN(n_2699));
   AOI21_X1 i_2438 (.A(n_3440), .B1(n_3439), .B2(n_2861), .ZN(n_2703));
   XNOR2_X1 i_2439 (.A(n_3605), .B(n_2709), .ZN(n_3607));
   INV_X1 i_2440 (.A(n_2709), .ZN(n_2704));
   AOI21_X1 i_2441 (.A(n_3430), .B1(n_3429), .B2(n_2858), .ZN(n_2709));
   INV_X1 i_2442 (.A(n_2713), .ZN(n_3448));
   AOI21_X1 i_2443 (.A(n_3445), .B1(n_3444), .B2(n_2865), .ZN(n_2713));
   XNOR2_X1 i_2444 (.A(n_3600), .B(n_2717), .ZN(n_3602));
   INV_X1 i_2445 (.A(n_2717), .ZN(n_2714));
   AOI21_X1 i_2446 (.A(n_3410), .B1(n_3409), .B2(n_2866), .ZN(n_2717));
   INV_X1 i_2447 (.A(n_2718), .ZN(n_3438));
   AOI21_X1 i_2448 (.A(n_3435), .B1(n_3434), .B2(n_2880), .ZN(n_2718));
   XOR2_X1 i_2449 (.A(n_3575), .B(n_2719), .Z(n_3577));
   XOR2_X1 i_2450 (.A(n_2721), .B(n_2720), .Z(n_2719));
   NAND2_X1 i_2451 (.A1(inputB[7]), .A2(inputA[24]), .ZN(n_2720));
   NAND2_X1 i_2452 (.A1(n_2725), .A2(n_2723), .ZN(n_2721));
   INV_X1 i_2453 (.A(n_2724), .ZN(n_2723));
   AOI22_X1 i_2454 (.A1(inputB[5]), .A2(inputA[26]), .B1(inputB[6]), .B2(
      inputA[25]), .ZN(n_2724));
   NAND3_X1 i_2455 (.A1(inputB[6]), .A2(inputA[26]), .A3(n_3013), .ZN(n_2725));
   XOR2_X1 i_2456 (.A(n_3580), .B(n_2726), .Z(n_3582));
   XOR2_X1 i_2457 (.A(n_2728), .B(n_2727), .Z(n_2726));
   NAND2_X1 i_2458 (.A1(inputB[16]), .A2(inputA[15]), .ZN(n_2727));
   NAND2_X1 i_2459 (.A1(n_2732), .A2(n_2729), .ZN(n_2728));
   INV_X1 i_2460 (.A(n_2731), .ZN(n_2729));
   AOI22_X1 i_2461 (.A1(inputB[14]), .A2(inputA[17]), .B1(inputB[15]), .B2(
      inputA[16]), .ZN(n_2731));
   NAND3_X1 i_2462 (.A1(inputB[15]), .A2(inputA[17]), .A3(n_2997), .ZN(n_2732));
   XNOR2_X1 i_2463 (.A(n_3590), .B(n_2734), .ZN(n_3592));
   INV_X1 i_2464 (.A(n_2734), .ZN(n_2733));
   AOI21_X1 i_2465 (.A(n_3400), .B1(n_3399), .B2(n_2923), .ZN(n_2734));
   INV_X1 i_2466 (.A(n_2735), .ZN(n_3428));
   AOI21_X1 i_2467 (.A(n_3425), .B1(n_3424), .B2(n_2878), .ZN(n_2735));
   XOR2_X1 i_2468 (.A(n_3570), .B(n_2738), .Z(n_3572));
   OAI21_X1 i_2469 (.A(n_2917), .B1(n_2916), .B2(n_2914), .ZN(n_2738));
   INV_X1 i_2470 (.A(n_2739), .ZN(n_3408));
   AOI21_X1 i_2471 (.A(n_3405), .B1(n_3404), .B2(n_2881), .ZN(n_2739));
   INV_X1 i_2472 (.A(n_2740), .ZN(n_3418));
   AOI21_X1 i_2473 (.A(n_3415), .B1(n_3414), .B2(n_2892), .ZN(n_2740));
   INV_X1 i_2474 (.A(n_2741), .ZN(n_3423));
   AOI21_X1 i_2475 (.A(n_3420), .B1(n_3419), .B2(n_2901), .ZN(n_2741));
   XOR2_X1 i_2476 (.A(n_3560), .B(n_2742), .Z(n_3562));
   AOI21_X1 i_2477 (.A(n_2896), .B1(n_2897), .B2(n_2893), .ZN(n_2742));
   XOR2_X1 i_2478 (.A(n_3565), .B(n_2744), .Z(n_3567));
   AOI22_X1 i_2479 (.A1(n_3106), .A2(n_2908), .B1(n_2906), .B2(n_2902), .ZN(
      n_2744));
   XNOR2_X1 i_2481 (.A(n_2747), .B(n_2746), .ZN(n_3477));
   INV_X1 i_2482 (.A(n_2746), .ZN(n_2745));
   NAND2_X1 i_2483 (.A1(inputB[31]), .A2(inputA[0]), .ZN(n_2746));
   NAND2_X1 i_2485 (.A1(n_2750), .A2(n_2748), .ZN(n_2747));
   OR2_X1 i_2486 (.A1(n_2908), .A2(n_2749), .ZN(n_2748));
   NAND2_X1 i_2487 (.A1(inputB[30]), .A2(inputA[2]), .ZN(n_2749));
   INV_X1 i_2489 (.A(n_2752), .ZN(n_2750));
   AOI22_X1 i_2490 (.A1(inputB[29]), .A2(inputA[2]), .B1(inputB[30]), .B2(
      inputA[1]), .ZN(n_2752));
   XOR2_X1 i_2491 (.A(n_2754), .B(n_2753), .Z(n_3486));
   NAND2_X1 i_2493 (.A1(inputB[28]), .A2(inputA[3]), .ZN(n_2753));
   NAND2_X1 i_2494 (.A1(n_2756), .A2(n_2755), .ZN(n_2754));
   NAND3_X1 i_2495 (.A1(inputB[26]), .A2(inputA[5]), .A3(n_2760), .ZN(n_2755));
   INV_X1 i_2497 (.A(n_2759), .ZN(n_2756));
   AOI21_X1 i_2498 (.A(n_2760), .B1(inputB[26]), .B2(inputA[5]), .ZN(n_2759));
   AND2_X1 i_2499 (.A1(inputB[27]), .A2(inputA[4]), .ZN(n_2760));
   XOR2_X1 i_2501 (.A(n_2762), .B(n_2761), .Z(n_3500));
   AND2_X1 i_2502 (.A1(inputB[22]), .A2(inputA[9]), .ZN(n_2761));
   AND2_X1 i_2503 (.A1(n_2765), .A2(n_2763), .ZN(n_2762));
   NAND2_X1 i_2505 (.A1(n_2900), .A2(n_2767), .ZN(n_2763));
   NAND2_X1 i_2506 (.A1(n_2899), .A2(n_2766), .ZN(n_2765));
   INV_X1 i_2507 (.A(n_2767), .ZN(n_2766));
   NAND2_X1 i_2509 (.A1(inputB[21]), .A2(inputA[10]), .ZN(n_2767));
   XOR2_X1 i_2510 (.A(n_2769), .B(n_2768), .Z(n_3507));
   NAND2_X1 i_2511 (.A1(inputB[19]), .A2(inputA[12]), .ZN(n_2768));
   NAND2_X1 i_2513 (.A1(n_2771), .A2(n_2770), .ZN(n_2769));
   NAND3_X1 i_2514 (.A1(inputB[17]), .A2(inputA[14]), .A3(n_2773), .ZN(n_2770));
   INV_X1 i_2515 (.A(n_2772), .ZN(n_2771));
   AOI21_X1 i_2517 (.A(n_2773), .B1(inputB[17]), .B2(inputA[14]), .ZN(n_2772));
   AND2_X1 i_2518 (.A1(inputB[18]), .A2(inputA[13]), .ZN(n_2773));
   XOR2_X1 i_2519 (.A(n_2775), .B(n_2774), .Z(n_3521));
   NAND2_X1 i_2521 (.A1(inputB[13]), .A2(inputA[18]), .ZN(n_2774));
   OAI21_X1 i_2522 (.A(n_2778), .B1(n_2871), .B2(n_2779), .ZN(n_2775));
   NAND2_X1 i_2523 (.A1(n_2871), .A2(n_2779), .ZN(n_2778));
   INV_X1 i_2525 (.A(n_2780), .ZN(n_2779));
   NAND2_X1 i_2526 (.A1(inputB[12]), .A2(inputA[19]), .ZN(n_2780));
   XOR2_X1 i_2527 (.A(n_2789), .B(n_2784), .Z(n_3528));
   NAND2_X1 i_2529 (.A1(inputB[10]), .A2(inputA[21]), .ZN(n_2784));
   NAND2_X1 i_2530 (.A1(n_2798), .A2(n_2794), .ZN(n_2789));
   NAND3_X1 i_2531 (.A1(inputB[8]), .A2(inputA[23]), .A3(n_2800), .ZN(n_2794));
   INV_X1 i_2533 (.A(n_2799), .ZN(n_2798));
   AOI21_X1 i_2534 (.A(n_2800), .B1(inputB[8]), .B2(inputA[23]), .ZN(n_2799));
   AND2_X1 i_2535 (.A1(inputB[9]), .A2(inputA[22]), .ZN(n_2800));
   XNOR2_X1 i_2537 (.A(n_2809), .B(n_2804), .ZN(n_3542));
   NAND2_X1 i_2538 (.A1(inputB[4]), .A2(inputA[27]), .ZN(n_2804));
   AND2_X1 i_2539 (.A1(n_2814), .A2(n_2813), .ZN(n_2809));
   NAND2_X1 i_2540 (.A1(n_2889), .A2(n_2819), .ZN(n_2813));
   OR2_X1 i_2541 (.A1(n_2889), .A2(n_2819), .ZN(n_2814));
   NAND2_X1 i_2542 (.A1(inputB[3]), .A2(inputA[28]), .ZN(n_2819));
   XNOR2_X1 i_2543 (.A(n_2825), .B(n_2824), .ZN(n_3549));
   OAI21_X1 i_2544 (.A(n_2888), .B1(n_2887), .B2(n_2882), .ZN(n_2824));
   NAND2_X1 i_2545 (.A1(n_2833), .A2(n_2829), .ZN(n_2825));
   INV_X1 i_2546 (.A(n_2830), .ZN(n_2829));
   AOI211_X1 i_2547 (.A(n_5754), .B(n_5751), .C1(inputB[0]), .C2(inputA[31]), 
      .ZN(n_2830));
   OAI211_X1 i_2548 (.A(inputB[0]), .B(inputA[31]), .C1(n_5754), .C2(n_5751), 
      .ZN(n_2833));
   INV_X1 i_2549 (.A(n_2834), .ZN(n_3393));
   AOI21_X1 i_2550 (.A(n_3390), .B1(n_3389), .B2(n_2922), .ZN(n_2834));
   INV_X1 i_2551 (.A(n_2835), .ZN(n_3398));
   AOI21_X1 i_2552 (.A(n_3395), .B1(n_3394), .B2(n_2879), .ZN(n_2835));
   OAI21_X1 i_2553 (.A(n_2936), .B1(n_2942), .B2(n_2932), .ZN(n_3321));
   OAI21_X1 i_2554 (.A(n_2951), .B1(n_2957), .B2(n_2947), .ZN(n_3328));
   OAI21_X1 i_2555 (.A(n_2972), .B1(n_2978), .B2(n_2963), .ZN(n_3342));
   OAI21_X1 i_2556 (.A(n_2992), .B1(n_2987), .B2(n_2981), .ZN(n_3349));
   OAI21_X1 i_2557 (.A(n_3003), .B1(n_3005), .B2(n_3001), .ZN(n_3363));
   OAI21_X1 i_2558 (.A(n_3008), .B1(n_3012), .B2(n_3006), .ZN(n_3370));
   XOR2_X1 i_2559 (.A(n_3469), .B(n_2839), .Z(n_3471));
   XNOR2_X1 i_2560 (.A(n_3464), .B(n_2844), .ZN(n_2839));
   INV_X1 i_2561 (.A(n_2844), .ZN(n_2843));
   AOI21_X1 i_2562 (.A(n_3295), .B1(n_3294), .B2(n_3024), .ZN(n_2844));
   INV_X1 i_2563 (.A(n_2849), .ZN(n_3308));
   AOI21_X1 i_2564 (.A(n_3305), .B1(n_3304), .B2(n_3020), .ZN(n_2849));
   XNOR2_X1 i_2565 (.A(n_3459), .B(n_2854), .ZN(n_3461));
   INV_X1 i_2566 (.A(n_2854), .ZN(n_2853));
   AOI21_X1 i_2567 (.A(n_3290), .B1(n_3289), .B2(n_3036), .ZN(n_2854));
   INV_X1 i_2568 (.A(n_2855), .ZN(n_3303));
   AOI21_X1 i_2569 (.A(n_3300), .B1(n_3299), .B2(n_3021), .ZN(n_2855));
   XOR2_X1 i_2570 (.A(n_3449), .B(n_2857), .Z(n_3451));
   XNOR2_X1 i_2571 (.A(n_3429), .B(n_2859), .ZN(n_2857));
   INV_X1 i_2572 (.A(n_2859), .ZN(n_2858));
   AOI21_X1 i_2573 (.A(n_3255), .B1(n_3254), .B2(n_3063), .ZN(n_2859));
   XOR2_X1 i_2574 (.A(n_3454), .B(n_2860), .Z(n_3456));
   XNOR2_X1 i_2575 (.A(n_3439), .B(n_2864), .ZN(n_2860));
   INV_X1 i_2576 (.A(n_2864), .ZN(n_2861));
   AOI21_X1 i_2577 (.A(n_3260), .B1(n_3259), .B2(n_3050), .ZN(n_2864));
   XOR2_X1 i_2578 (.A(n_3444), .B(n_2865), .Z(n_3446));
   XOR2_X1 i_2579 (.A(n_3409), .B(n_2866), .Z(n_2865));
   XOR2_X1 i_2580 (.A(n_2868), .B(n_2867), .Z(n_2866));
   NAND2_X1 i_2581 (.A1(inputB[12]), .A2(inputA[18]), .ZN(n_2867));
   NAND2_X1 i_2582 (.A1(n_2873), .A2(n_2870), .ZN(n_2868));
   NAND2_X1 i_2583 (.A1(n_3163), .A2(n_2871), .ZN(n_2870));
   INV_X1 i_2584 (.A(n_2872), .ZN(n_2871));
   NAND2_X1 i_2585 (.A1(inputB[11]), .A2(inputA[20]), .ZN(n_2872));
   INV_X1 i_2586 (.A(n_2874), .ZN(n_2873));
   AOI22_X1 i_2587 (.A1(inputB[10]), .A2(inputA[20]), .B1(inputB[11]), .B2(
      inputA[19]), .ZN(n_2874));
   INV_X1 i_2588 (.A(n_2875), .ZN(n_3288));
   AOI21_X1 i_2589 (.A(n_3285), .B1(n_3284), .B2(n_3041), .ZN(n_2875));
   INV_X1 i_2590 (.A(n_2876), .ZN(n_3283));
   AOI21_X1 i_2591 (.A(n_3280), .B1(n_3279), .B2(n_3025), .ZN(n_2876));
   XOR2_X1 i_2592 (.A(n_3424), .B(n_2878), .Z(n_3426));
   XOR2_X1 i_2593 (.A(n_3394), .B(n_2879), .Z(n_2878));
   OAI21_X1 i_2594 (.A(n_3120), .B1(n_3125), .B2(n_3114), .ZN(n_2879));
   XOR2_X1 i_2595 (.A(n_3434), .B(n_2880), .Z(n_3436));
   XOR2_X1 i_2596 (.A(n_3404), .B(n_2881), .Z(n_2880));
   XOR2_X1 i_2597 (.A(n_2885), .B(n_2882), .Z(n_2881));
   NAND2_X1 i_2598 (.A1(inputB[3]), .A2(inputA[27]), .ZN(n_2882));
   NAND2_X1 i_2599 (.A1(n_2888), .A2(n_2886), .ZN(n_2885));
   INV_X1 i_2601 (.A(n_2887), .ZN(n_2886));
   AOI22_X1 i_2602 (.A1(inputB[1]), .A2(inputA[29]), .B1(inputB[2]), .B2(
      inputA[28]), .ZN(n_2887));
   NAND3_X1 i_2603 (.A1(inputB[2]), .A2(inputA[29]), .A3(n_3258), .ZN(n_2888));
   NAND2_X1 i_2605 (.A1(inputB[2]), .A2(inputA[29]), .ZN(n_2889));
   INV_X1 i_2606 (.A(n_2891), .ZN(n_3278));
   AOI21_X1 i_2607 (.A(n_3275), .B1(n_3274), .B2(n_3037), .ZN(n_2891));
   XOR2_X1 i_2609 (.A(n_3414), .B(n_2892), .Z(n_3416));
   XOR2_X1 i_2610 (.A(n_2894), .B(n_2893), .Z(n_2892));
   NAND2_X1 i_2611 (.A1(inputB[21]), .A2(inputA[9]), .ZN(n_2893));
   NAND2_X1 i_2613 (.A1(n_2897), .A2(n_2895), .ZN(n_2894));
   INV_X1 i_2614 (.A(n_2896), .ZN(n_2895));
   AOI22_X1 i_2615 (.A1(inputB[19]), .A2(inputA[11]), .B1(inputB[20]), .B2(
      inputA[10]), .ZN(n_2896));
   NAND2_X1 i_2617 (.A1(n_3141), .A2(n_2899), .ZN(n_2897));
   INV_X1 i_2618 (.A(n_2900), .ZN(n_2899));
   NAND2_X1 i_2619 (.A1(inputB[20]), .A2(inputA[11]), .ZN(n_2900));
   XOR2_X1 i_2621 (.A(n_3419), .B(n_2901), .Z(n_3421));
   XOR2_X1 i_2622 (.A(n_2903), .B(n_2902), .Z(n_2901));
   NAND2_X1 i_2623 (.A1(inputB[30]), .A2(inputA[0]), .ZN(n_2902));
   OAI21_X1 i_2625 (.A(n_2906), .B1(n_3105), .B2(n_2907), .ZN(n_2903));
   NAND2_X1 i_2626 (.A1(n_3105), .A2(n_2907), .ZN(n_2906));
   INV_X1 i_2627 (.A(n_2908), .ZN(n_2907));
   NAND2_X1 i_2629 (.A1(inputB[29]), .A2(inputA[1]), .ZN(n_2908));
   INV_X1 i_2630 (.A(n_2909), .ZN(n_3268));
   AOI21_X1 i_2631 (.A(n_3265), .B1(n_3264), .B2(n_3047), .ZN(n_2909));
   INV_X1 i_2633 (.A(n_2910), .ZN(n_3273));
   AOI21_X1 i_2634 (.A(n_3270), .B1(n_3269), .B2(n_3042), .ZN(n_2910));
   INV_X1 i_2635 (.A(n_2912), .ZN(n_3248));
   AOI21_X1 i_2637 (.A(n_3245), .B1(n_3244), .B2(n_3026), .ZN(n_2912));
   INV_X1 i_2638 (.A(n_2913), .ZN(n_3253));
   AOI21_X1 i_2639 (.A(n_3250), .B1(n_3249), .B2(n_3054), .ZN(n_2913));
   XNOR2_X1 i_2641 (.A(n_2915), .B(n_2914), .ZN(n_3383));
   NAND2_X1 i_2642 (.A1(inputB[0]), .A2(inputA[30]), .ZN(n_2914));
   AOI21_X1 i_2643 (.A(n_2916), .B1(n_2921), .B2(n_2920), .ZN(n_2915));
   NOR2_X1 i_2645 (.A1(n_2921), .A2(n_2920), .ZN(n_2916));
   NAND2_X1 i_2646 (.A1(n_2921), .A2(n_2920), .ZN(n_2917));
   OAI21_X1 i_2647 (.A(n_3168), .B1(n_3171), .B2(n_3166), .ZN(n_2920));
   OAI21_X1 i_2649 (.A(n_3174), .B1(n_3176), .B2(n_3172), .ZN(n_2921));
   XOR2_X1 i_2650 (.A(n_3389), .B(n_2922), .Z(n_3391));
   OAI21_X1 i_2651 (.A(n_3154), .B1(n_3158), .B2(n_3145), .ZN(n_2922));
   XNOR2_X1 i_2653 (.A(n_3399), .B(n_2926), .ZN(n_3401));
   INV_X1 i_2654 (.A(n_2926), .ZN(n_2923));
   AOI21_X1 i_2655 (.A(n_3235), .B1(n_3234), .B2(n_3051), .ZN(n_2926));
   INV_X1 i_2657 (.A(n_2927), .ZN(n_3243));
   AOI21_X1 i_2658 (.A(n_3240), .B1(n_3239), .B2(n_3071), .ZN(n_2927));
   XOR2_X1 i_2659 (.A(n_2933), .B(n_2932), .Z(n_3320));
   NAND2_X1 i_2661 (.A1(inputB[27]), .A2(inputA[3]), .ZN(n_2932));
   NAND2_X1 i_2662 (.A1(n_2937), .A2(n_2936), .ZN(n_2933));
   NAND3_X1 i_2663 (.A1(inputB[26]), .A2(inputA[4]), .A3(n_3069), .ZN(n_2936));
   INV_X1 i_2664 (.A(n_2942), .ZN(n_2937));
   AOI21_X1 i_2665 (.A(n_3069), .B1(inputB[26]), .B2(inputA[4]), .ZN(n_2942));
   XOR2_X1 i_2666 (.A(n_2948), .B(n_2947), .Z(n_3327));
   NAND2_X1 i_2667 (.A1(inputB[24]), .A2(inputA[6]), .ZN(n_2947));
   NAND2_X1 i_2668 (.A1(n_2952), .A2(n_2951), .ZN(n_2948));
   NAND3_X1 i_2669 (.A1(inputB[22]), .A2(inputA[8]), .A3(n_2962), .ZN(n_2951));
   INV_X1 i_2670 (.A(n_2957), .ZN(n_2952));
   AOI21_X1 i_2671 (.A(n_2962), .B1(inputB[22]), .B2(inputA[8]), .ZN(n_2957));
   AND2_X1 i_2672 (.A1(inputB[23]), .A2(inputA[7]), .ZN(n_2962));
   XOR2_X1 i_2673 (.A(n_2967), .B(n_2963), .Z(n_3341));
   NAND2_X1 i_2674 (.A1(inputB[18]), .A2(inputA[12]), .ZN(n_2963));
   NAND2_X1 i_2675 (.A1(n_2977), .A2(n_2972), .ZN(n_2967));
   NAND3_X1 i_2676 (.A1(inputB[17]), .A2(inputA[13]), .A3(n_3062), .ZN(n_2972));
   INV_X1 i_2677 (.A(n_2978), .ZN(n_2977));
   AOI21_X1 i_2678 (.A(n_3062), .B1(inputB[17]), .B2(inputA[13]), .ZN(n_2978));
   XNOR2_X1 i_2679 (.A(n_2982), .B(n_2981), .ZN(n_3348));
   NAND2_X1 i_2680 (.A1(inputB[15]), .A2(inputA[15]), .ZN(n_2981));
   NOR2_X1 i_2681 (.A1(n_2991), .A2(n_2987), .ZN(n_2982));
   AOI21_X1 i_2682 (.A(n_2997), .B1(inputB[13]), .B2(inputA[17]), .ZN(n_2987));
   INV_X1 i_2683 (.A(n_2992), .ZN(n_2991));
   NAND3_X1 i_2684 (.A1(inputB[13]), .A2(inputA[17]), .A3(n_2997), .ZN(n_2992));
   AND2_X1 i_2685 (.A1(inputB[14]), .A2(inputA[16]), .ZN(n_2997));
   XOR2_X1 i_2686 (.A(n_3002), .B(n_3001), .Z(n_3362));
   NAND2_X1 i_2687 (.A1(inputB[9]), .A2(inputA[21]), .ZN(n_3001));
   NAND2_X1 i_2688 (.A1(n_3004), .A2(n_3003), .ZN(n_3002));
   NAND3_X1 i_2689 (.A1(inputB[8]), .A2(inputA[22]), .A3(n_3034), .ZN(n_3003));
   INV_X1 i_2690 (.A(n_3005), .ZN(n_3004));
   AOI21_X1 i_2691 (.A(n_3034), .B1(inputB[8]), .B2(inputA[22]), .ZN(n_3005));
   XOR2_X1 i_2692 (.A(n_3007), .B(n_3006), .Z(n_3369));
   NAND2_X1 i_2693 (.A1(inputB[6]), .A2(inputA[24]), .ZN(n_3006));
   NAND2_X1 i_2694 (.A1(n_3009), .A2(n_3008), .ZN(n_3007));
   NAND3_X1 i_2695 (.A1(inputB[4]), .A2(inputA[26]), .A3(n_3013), .ZN(n_3008));
   INV_X1 i_2696 (.A(n_3012), .ZN(n_3009));
   AOI21_X1 i_2697 (.A(n_3013), .B1(inputB[4]), .B2(inputA[26]), .ZN(n_3012));
   AND2_X1 i_2698 (.A1(inputB[5]), .A2(inputA[25]), .ZN(n_3013));
   INV_X1 i_2699 (.A(n_3014), .ZN(n_3228));
   AOI21_X1 i_2700 (.A(n_3225), .B1(n_3224), .B2(n_3085), .ZN(n_3014));
   INV_X1 i_2701 (.A(n_3015), .ZN(n_3233));
   AOI21_X1 i_2702 (.A(n_3230), .B1(n_3229), .B2(n_3090), .ZN(n_3015));
   OAI21_X1 i_2703 (.A(n_3100), .B1(n_3111), .B2(n_3095), .ZN(n_3157));
   OAI21_X1 i_2704 (.A(n_3068), .B1(n_3067), .B2(n_3064), .ZN(n_3164));
   NAND2_X1 i_2705 (.A1(n_3140), .A2(n_3016), .ZN(n_3178));
   NAND2_X1 i_2706 (.A1(n_3135), .A2(n_3130), .ZN(n_3016));
   OAI21_X1 i_2707 (.A(n_3061), .B1(n_3058), .B2(n_3055), .ZN(n_3185));
   NAND2_X1 i_2708 (.A1(n_3162), .A2(n_3019), .ZN(n_3199));
   NAND2_X1 i_2709 (.A1(n_3161), .A2(n_3159), .ZN(n_3019));
   OAI21_X1 i_2710 (.A(n_3033), .B1(n_3030), .B2(n_3027), .ZN(n_3206));
   XOR2_X1 i_2711 (.A(n_3304), .B(n_3020), .Z(n_3306));
   XNOR2_X1 i_2712 (.A(n_3299), .B(n_3022), .ZN(n_3020));
   INV_X1 i_2713 (.A(n_3022), .ZN(n_3021));
   AOI21_X1 i_2714 (.A(n_3138), .B1(n_3137), .B2(n_3188), .ZN(n_3022));
   INV_X1 i_2715 (.A(n_3023), .ZN(n_3151));
   AOI21_X1 i_2716 (.A(n_3148), .B1(n_3147), .B2(n_3181), .ZN(n_3023));
   XOR2_X1 i_2717 (.A(n_3294), .B(n_3024), .Z(n_3296));
   XOR2_X1 i_2718 (.A(n_3279), .B(n_3025), .Z(n_3024));
   XOR2_X1 i_2719 (.A(n_3244), .B(n_3026), .Z(n_3025));
   XOR2_X1 i_2720 (.A(n_3028), .B(n_3027), .Z(n_3026));
   NAND2_X1 i_2721 (.A1(inputB[8]), .A2(inputA[21]), .ZN(n_3027));
   NAND2_X1 i_2722 (.A1(n_3033), .A2(n_3029), .ZN(n_3028));
   INV_X1 i_2723 (.A(n_3030), .ZN(n_3029));
   AOI22_X1 i_2724 (.A1(inputB[6]), .A2(inputA[23]), .B1(inputB[7]), .B2(
      inputA[22]), .ZN(n_3030));
   NAND2_X1 i_2725 (.A1(n_3330), .A2(n_3034), .ZN(n_3033));
   AND2_X1 i_2726 (.A1(inputB[7]), .A2(inputA[23]), .ZN(n_3034));
   INV_X1 i_2727 (.A(n_3035), .ZN(n_3146));
   AOI21_X1 i_2728 (.A(n_3143), .B1(n_3142), .B2(n_3182), .ZN(n_3035));
   XOR2_X1 i_2729 (.A(n_3289), .B(n_3036), .Z(n_3291));
   XNOR2_X1 i_2730 (.A(n_3274), .B(n_3040), .ZN(n_3036));
   INV_X1 i_2731 (.A(n_3040), .ZN(n_3037));
   AOI21_X1 i_2733 (.A(n_3108), .B1(n_3107), .B2(n_3210), .ZN(n_3040));
   XOR2_X1 i_2734 (.A(n_3284), .B(n_3041), .Z(n_3286));
   XNOR2_X1 i_2735 (.A(n_3269), .B(n_3043), .ZN(n_3041));
   INV_X1 i_2737 (.A(n_3043), .ZN(n_3042));
   AOI21_X1 i_2738 (.A(n_3088), .B1(n_3087), .B2(n_3246), .ZN(n_3043));
   INV_X1 i_2739 (.A(n_3044), .ZN(n_3136));
   AOI21_X1 i_2741 (.A(n_3133), .B1(n_3132), .B2(n_3183), .ZN(n_3044));
   INV_X1 i_2742 (.A(n_3045), .ZN(n_3131));
   AOI21_X1 i_2743 (.A(n_3128), .B1(n_3127), .B2(n_3202), .ZN(n_3045));
   INV_X1 i_2745 (.A(n_3046), .ZN(n_3126));
   AOI21_X1 i_2746 (.A(n_3123), .B1(n_3122), .B2(n_3189), .ZN(n_3046));
   XNOR2_X1 i_2747 (.A(n_3264), .B(n_3048), .ZN(n_3266));
   INV_X1 i_2749 (.A(n_3048), .ZN(n_3047));
   AOI21_X1 i_2750 (.A(n_3103), .B1(n_3102), .B2(n_3223), .ZN(n_3048));
   INV_X1 i_2751 (.A(n_3049), .ZN(n_3121));
   AOI21_X1 i_2753 (.A(n_3118), .B1(n_3117), .B2(n_3207), .ZN(n_3049));
   XOR2_X1 i_2754 (.A(n_3259), .B(n_3050), .Z(n_3261));
   XOR2_X1 i_2755 (.A(n_3234), .B(n_3051), .Z(n_3050));
   AOI22_X1 i_2757 (.A1(n_3364), .A2(n_3238), .B1(n_3236), .B2(n_3227), .ZN(
      n_3051));
   XOR2_X1 i_2758 (.A(n_3249), .B(n_3054), .Z(n_3251));
   XOR2_X1 i_2759 (.A(n_3056), .B(n_3055), .Z(n_3054));
   NAND2_X1 i_2761 (.A1(inputB[17]), .A2(inputA[12]), .ZN(n_3055));
   NAND2_X1 i_2762 (.A1(n_3061), .A2(n_3057), .ZN(n_3056));
   INV_X1 i_2763 (.A(n_3058), .ZN(n_3057));
   AOI22_X1 i_2765 (.A1(inputB[15]), .A2(inputA[14]), .B1(inputB[16]), .B2(
      inputA[13]), .ZN(n_3058));
   NAND2_X1 i_2766 (.A1(n_3315), .A2(n_3062), .ZN(n_3061));
   AND2_X1 i_2767 (.A1(inputB[16]), .A2(inputA[14]), .ZN(n_3062));
   XOR2_X1 i_2769 (.A(n_3254), .B(n_3063), .Z(n_3256));
   XOR2_X1 i_2770 (.A(n_3065), .B(n_3064), .Z(n_3063));
   NAND2_X1 i_2771 (.A1(inputB[26]), .A2(inputA[3]), .ZN(n_3064));
   NAND2_X1 i_2773 (.A1(n_3068), .A2(n_3066), .ZN(n_3065));
   INV_X1 i_2774 (.A(n_3067), .ZN(n_3066));
   AOI22_X1 i_2775 (.A1(inputB[24]), .A2(inputA[5]), .B1(inputB[25]), .B2(
      inputA[4]), .ZN(n_3067));
   NAND2_X1 i_2777 (.A1(n_3293), .A2(n_3069), .ZN(n_3068));
   AND2_X1 i_2778 (.A1(inputB[25]), .A2(inputA[5]), .ZN(n_3069));
   INV_X1 i_2779 (.A(n_3070), .ZN(n_3116));
   AOI21_X1 i_2781 (.A(n_3113), .B1(n_3112), .B2(n_3203), .ZN(n_3070));
   XNOR2_X1 i_2782 (.A(n_3239), .B(n_3075), .ZN(n_3241));
   INV_X1 i_2783 (.A(n_3075), .ZN(n_3071));
   AOI22_X1 i_2785 (.A1(n_3403), .A2(n_3258), .B1(n_3252), .B2(n_3247), .ZN(
      n_3075));
   INV_X1 i_2786 (.A(n_3079), .ZN(n_3096));
   AOI21_X1 i_2787 (.A(n_3093), .B1(n_3092), .B2(n_3214), .ZN(n_3079));
   INV_X1 i_2789 (.A(n_3080), .ZN(n_3101));
   AOI21_X1 i_2790 (.A(n_3098), .B1(n_3097), .B2(n_3190), .ZN(n_3080));
   XOR2_X1 i_2791 (.A(n_3224), .B(n_3085), .Z(n_3226));
   AOI21_X1 i_2793 (.A(n_3217), .B1(n_3220), .B2(n_3215), .ZN(n_3085));
   XOR2_X1 i_2794 (.A(n_3229), .B(n_3090), .Z(n_3231));
   AOI21_X1 i_2795 (.A(n_3200), .B1(n_3195), .B2(n_3192), .ZN(n_3090));
   INV_X1 i_2796 (.A(n_3091), .ZN(n_3086));
   AOI21_X1 i_2797 (.A(n_3083), .B1(n_3082), .B2(n_3271), .ZN(n_3091));
   XOR2_X1 i_2798 (.A(n_3099), .B(n_3095), .Z(n_3156));
   NAND2_X1 i_2799 (.A1(inputB[29]), .A2(inputA[0]), .ZN(n_3095));
   NAND2_X1 i_2800 (.A1(n_3110), .A2(n_3100), .ZN(n_3099));
   NAND2_X1 i_2801 (.A1(n_3237), .A2(n_3105), .ZN(n_3100));
   INV_X1 i_2802 (.A(n_3106), .ZN(n_3105));
   NAND2_X1 i_2803 (.A1(inputB[28]), .A2(inputA[2]), .ZN(n_3106));
   INV_X1 i_2804 (.A(n_3111), .ZN(n_3110));
   AOI22_X1 i_2805 (.A1(inputB[27]), .A2(inputA[2]), .B1(inputB[28]), .B2(
      inputA[1]), .ZN(n_3111));
   XOR2_X1 i_2806 (.A(n_3115), .B(n_3114), .Z(n_3170));
   NAND2_X1 i_2807 (.A1(inputB[23]), .A2(inputA[6]), .ZN(n_3114));
   NAND2_X1 i_2808 (.A1(n_3124), .A2(n_3120), .ZN(n_3115));
   NAND3_X1 i_2809 (.A1(inputB[22]), .A2(inputA[7]), .A3(n_3302), .ZN(n_3120));
   INV_X1 i_2810 (.A(n_3125), .ZN(n_3124));
   AOI21_X1 i_2811 (.A(n_3302), .B1(inputB[22]), .B2(inputA[7]), .ZN(n_3125));
   XOR2_X1 i_2812 (.A(n_3134), .B(n_3130), .Z(n_3177));
   AND2_X1 i_2813 (.A1(inputB[20]), .A2(inputA[9]), .ZN(n_3130));
   AND2_X1 i_2814 (.A1(n_3140), .A2(n_3135), .ZN(n_3134));
   NAND2_X1 i_2815 (.A1(n_3197), .A2(n_3144), .ZN(n_3135));
   NAND2_X1 i_2816 (.A1(n_3196), .A2(n_3141), .ZN(n_3140));
   INV_X1 i_2817 (.A(n_3144), .ZN(n_3141));
   NAND2_X1 i_2818 (.A1(inputB[19]), .A2(inputA[10]), .ZN(n_3144));
   XOR2_X1 i_2819 (.A(n_3150), .B(n_3145), .Z(n_3191));
   NAND2_X1 i_2820 (.A1(inputB[14]), .A2(inputA[15]), .ZN(n_3145));
   NAND2_X1 i_2821 (.A1(n_3155), .A2(n_3154), .ZN(n_3150));
   NAND3_X1 i_2822 (.A1(inputB[13]), .A2(inputA[16]), .A3(n_3322), .ZN(n_3154));
   INV_X1 i_2823 (.A(n_3158), .ZN(n_3155));
   AOI21_X1 i_2824 (.A(n_3322), .B1(inputB[13]), .B2(inputA[16]), .ZN(n_3158));
   XOR2_X1 i_2825 (.A(n_3160), .B(n_3159), .Z(n_3198));
   AND2_X1 i_2826 (.A1(inputB[11]), .A2(inputA[18]), .ZN(n_3159));
   AND2_X1 i_2827 (.A1(n_3162), .A2(n_3161), .ZN(n_3160));
   NAND2_X1 i_2828 (.A1(n_3222), .A2(n_3165), .ZN(n_3161));
   NAND2_X1 i_2829 (.A1(n_3221), .A2(n_3163), .ZN(n_3162));
   INV_X1 i_2830 (.A(n_3165), .ZN(n_3163));
   NAND2_X1 i_2831 (.A1(inputB[10]), .A2(inputA[19]), .ZN(n_3165));
   XOR2_X1 i_2832 (.A(n_3167), .B(n_3166), .Z(n_3212));
   NAND2_X1 i_2833 (.A1(inputB[5]), .A2(inputA[24]), .ZN(n_3166));
   NAND2_X1 i_2834 (.A1(n_3169), .A2(n_3168), .ZN(n_3167));
   NAND4_X1 i_2835 (.A1(inputB[3]), .A2(inputA[26]), .A3(inputB[4]), .A4(
      inputA[25]), .ZN(n_3168));
   INV_X1 i_2836 (.A(n_3171), .ZN(n_3169));
   AOI22_X1 i_2837 (.A1(inputB[3]), .A2(inputA[26]), .B1(inputB[4]), .B2(
      inputA[25]), .ZN(n_3171));
   XOR2_X1 i_2838 (.A(n_3173), .B(n_3172), .Z(n_3219));
   NAND2_X1 i_2839 (.A1(inputB[2]), .A2(inputA[27]), .ZN(n_3172));
   NAND2_X1 i_2840 (.A1(n_3175), .A2(n_3174), .ZN(n_3173));
   NAND3_X1 i_2841 (.A1(inputB[0]), .A2(inputA[29]), .A3(n_3258), .ZN(n_3174));
   INV_X1 i_2842 (.A(n_3176), .ZN(n_3175));
   AOI21_X1 i_2843 (.A(n_3258), .B1(inputB[0]), .B2(inputA[29]), .ZN(n_3176));
   INV_X1 i_2844 (.A(n_3179), .ZN(n_3076));
   AOI21_X1 i_2845 (.A(n_3073), .B1(n_3072), .B2(n_3267), .ZN(n_3179));
   INV_X1 i_2846 (.A(n_3180), .ZN(n_3081));
   AOI21_X1 i_2847 (.A(n_3078), .B1(n_3077), .B2(n_3211), .ZN(n_3180));
   OAI21_X1 i_2848 (.A(n_3282), .B1(n_3292), .B2(n_3277), .ZN(n_3011));
   OAI21_X1 i_2849 (.A(n_3301), .B1(n_3311), .B2(n_3297), .ZN(n_3018));
   AOI22_X1 i_2850 (.A1(n_3466), .A2(n_3316), .B1(n_3314), .B2(n_3312), .ZN(
      n_3032));
   OAI21_X1 i_2851 (.A(n_3319), .B1(n_3324), .B2(n_3317), .ZN(n_3039));
   AOI22_X1 i_2852 (.A1(n_3488), .A2(n_3331), .B1(n_3329), .B2(n_3325), .ZN(
      n_3053));
   OAI21_X1 i_2853 (.A(n_3336), .B1(n_3334), .B2(n_3332), .ZN(n_3060));
   XOR2_X1 i_2854 (.A(n_3147), .B(n_3181), .Z(n_3149));
   XOR2_X1 i_2855 (.A(n_3142), .B(n_3182), .Z(n_3181));
   XNOR2_X1 i_2856 (.A(n_3132), .B(n_3184), .ZN(n_3182));
   INV_X1 i_2857 (.A(n_3184), .ZN(n_3183));
   AOI21_X1 i_2858 (.A(n_2975), .B1(n_2974), .B2(n_3352), .ZN(n_3184));
   INV_X1 i_2859 (.A(n_3186), .ZN(n_2998));
   AOI21_X1 i_2860 (.A(n_2995), .B1(n_2994), .B2(n_3339), .ZN(n_3186));
   INV_X1 i_2861 (.A(n_3187), .ZN(n_2993));
   AOI21_X1 i_2862 (.A(n_2990), .B1(n_2989), .B2(n_3340), .ZN(n_3187));
   XOR2_X1 i_2863 (.A(n_3137), .B(n_3188), .Z(n_3139));
   XOR2_X1 i_2865 (.A(n_3122), .B(n_3189), .Z(n_3188));
   XOR2_X1 i_2866 (.A(n_3097), .B(n_3190), .Z(n_3189));
   XNOR2_X1 i_2867 (.A(n_3193), .B(n_3192), .ZN(n_3190));
   NAND2_X1 i_2869 (.A1(inputB[19]), .A2(inputA[9]), .ZN(n_3192));
   NOR2_X1 i_2870 (.A1(n_3200), .A2(n_3194), .ZN(n_3193));
   INV_X1 i_2871 (.A(n_3195), .ZN(n_3194));
   NAND3_X1 i_2873 (.A1(inputB[17]), .A2(inputA[10]), .A3(n_3196), .ZN(n_3195));
   INV_X1 i_2874 (.A(n_3197), .ZN(n_3196));
   NAND2_X1 i_2875 (.A1(inputB[18]), .A2(inputA[11]), .ZN(n_3197));
   AOI22_X1 i_2877 (.A1(inputB[17]), .A2(inputA[11]), .B1(inputB[18]), .B2(
      inputA[10]), .ZN(n_3200));
   INV_X1 i_2878 (.A(n_3201), .ZN(n_2988));
   AOI21_X1 i_2879 (.A(n_2985), .B1(n_2984), .B2(n_3347), .ZN(n_3201));
   XOR2_X1 i_2881 (.A(n_3127), .B(n_3202), .Z(n_3129));
   XNOR2_X1 i_2882 (.A(n_3112), .B(n_3204), .ZN(n_3202));
   INV_X1 i_2883 (.A(n_3204), .ZN(n_3203));
   AOI21_X1 i_2885 (.A(n_2945), .B1(n_2944), .B2(n_3381), .ZN(n_3204));
   INV_X1 i_2886 (.A(n_3205), .ZN(n_2983));
   AOI21_X1 i_2887 (.A(n_2980), .B1(n_2979), .B2(n_3343), .ZN(n_3205));
   XNOR2_X1 i_2889 (.A(n_3117), .B(n_3208), .ZN(n_3119));
   INV_X1 i_2890 (.A(n_3208), .ZN(n_3207));
   AOI21_X1 i_2891 (.A(n_2960), .B1(n_2959), .B2(n_3373), .ZN(n_3208));
   INV_X1 i_2893 (.A(n_3209), .ZN(n_2973));
   AOI21_X1 i_2894 (.A(n_2970), .B1(n_2969), .B2(n_3354), .ZN(n_3209));
   XOR2_X1 i_2895 (.A(n_3107), .B(n_3210), .Z(n_3109));
   XOR2_X1 i_2897 (.A(n_3077), .B(n_3211), .Z(n_3210));
   AOI22_X1 i_2898 (.A1(n_3545), .A2(n_3452), .B1(n_3443), .B2(n_3441), .ZN(
      n_3211));
   INV_X1 i_2899 (.A(n_3213), .ZN(n_2968));
   AOI21_X1 i_2901 (.A(n_2965), .B1(n_2964), .B2(n_3365), .ZN(n_3213));
   XOR2_X1 i_2902 (.A(n_3092), .B(n_3214), .Z(n_3094));
   XNOR2_X1 i_2903 (.A(n_3216), .B(n_3215), .ZN(n_3214));
   NAND2_X1 i_2905 (.A1(inputB[10]), .A2(inputA[18]), .ZN(n_3215));
   NOR2_X1 i_2906 (.A1(n_3218), .A2(n_3217), .ZN(n_3216));
   AOI22_X1 i_2907 (.A1(inputB[8]), .A2(inputA[20]), .B1(inputB[9]), .B2(
      inputA[19]), .ZN(n_3217));
   INV_X1 i_2909 (.A(n_3220), .ZN(n_3218));
   NAND3_X1 i_2910 (.A1(inputB[8]), .A2(inputA[19]), .A3(n_3221), .ZN(n_3220));
   INV_X1 i_2911 (.A(n_3222), .ZN(n_3221));
   NAND2_X1 i_2913 (.A1(inputB[9]), .A2(inputA[20]), .ZN(n_3222));
   XOR2_X1 i_2914 (.A(n_3102), .B(n_3223), .Z(n_3104));
   XOR2_X1 i_2915 (.A(n_3232), .B(n_3227), .Z(n_3223));
   NAND2_X1 i_2917 (.A1(inputB[28]), .A2(inputA[0]), .ZN(n_3227));
   OAI21_X1 i_2918 (.A(n_3236), .B1(n_3361), .B2(n_3237), .ZN(n_3232));
   NAND2_X1 i_2919 (.A1(n_3361), .A2(n_3237), .ZN(n_3236));
   INV_X1 i_2921 (.A(n_3238), .ZN(n_3237));
   NAND2_X1 i_2922 (.A1(inputB[27]), .A2(inputA[1]), .ZN(n_3238));
   INV_X1 i_2923 (.A(n_3242), .ZN(n_2958));
   AOI21_X1 i_2925 (.A(n_2955), .B1(n_2954), .B2(n_3368), .ZN(n_3242));
   XOR2_X1 i_2926 (.A(n_3087), .B(n_3246), .Z(n_3089));
   XOR2_X1 i_2927 (.A(n_3252), .B(n_3247), .Z(n_3246));
   OAI21_X1 i_2929 (.A(n_3496), .B1(n_3495), .B2(n_3491), .ZN(n_3247));
   AOI21_X1 i_2930 (.A(n_3257), .B1(n_3403), .B2(n_3258), .ZN(n_3252));
   AOI22_X1 i_2931 (.A1(inputB[0]), .A2(inputA[28]), .B1(inputB[1]), .B2(
      inputA[27]), .ZN(n_3257));
   AND2_X1 i_2932 (.A1(inputB[1]), .A2(inputA[28]), .ZN(n_3258));
   INV_X1 i_2933 (.A(n_3262), .ZN(n_2943));
   AOI21_X1 i_2934 (.A(n_2940), .B1(n_2939), .B2(n_3375), .ZN(n_3262));
   INV_X1 i_2935 (.A(n_3263), .ZN(n_2953));
   AOI21_X1 i_2936 (.A(n_2950), .B1(n_2949), .B2(n_3355), .ZN(n_3263));
   XOR2_X1 i_2937 (.A(n_3072), .B(n_3267), .Z(n_3074));
   AOI22_X1 i_2938 (.A1(n_3526), .A2(n_3481), .B1(n_3479), .B2(n_3476), .ZN(
      n_3267));
   XNOR2_X1 i_2939 (.A(n_3082), .B(n_3272), .ZN(n_3084));
   INV_X1 i_2940 (.A(n_3272), .ZN(n_3271));
   AOI21_X1 i_2941 (.A(n_2930), .B1(n_2929), .B2(n_3417), .ZN(n_3272));
   INV_X1 i_2942 (.A(n_3276), .ZN(n_2938));
   AOI21_X1 i_2943 (.A(n_2935), .B1(n_2934), .B2(n_3366), .ZN(n_3276));
   XOR2_X1 i_2944 (.A(n_3281), .B(n_3277), .Z(n_3010));
   NAND2_X1 i_2945 (.A1(inputB[25]), .A2(inputA[3]), .ZN(n_3277));
   NAND2_X1 i_2946 (.A1(n_3287), .A2(n_3282), .ZN(n_3281));
   NAND3_X1 i_2947 (.A1(inputB[23]), .A2(inputA[5]), .A3(n_3293), .ZN(n_3282));
   INV_X1 i_2948 (.A(n_3292), .ZN(n_3287));
   AOI21_X1 i_2949 (.A(n_3293), .B1(inputB[23]), .B2(inputA[5]), .ZN(n_3292));
   AND2_X1 i_2950 (.A1(inputB[24]), .A2(inputA[4]), .ZN(n_3293));
   XOR2_X1 i_2951 (.A(n_3298), .B(n_3297), .Z(n_3017));
   NAND2_X1 i_2952 (.A1(inputB[22]), .A2(inputA[6]), .ZN(n_3297));
   NAND2_X1 i_2953 (.A1(n_3307), .A2(n_3301), .ZN(n_3298));
   NAND2_X1 i_2954 (.A1(n_3447), .A2(n_3302), .ZN(n_3301));
   AND2_X1 i_2955 (.A1(inputB[21]), .A2(inputA[8]), .ZN(n_3302));
   INV_X1 i_2956 (.A(n_3311), .ZN(n_3307));
   AOI22_X1 i_2957 (.A1(inputB[20]), .A2(inputA[8]), .B1(inputB[21]), .B2(
      inputA[7]), .ZN(n_3311));
   XOR2_X1 i_2958 (.A(n_3313), .B(n_3312), .Z(n_3031));
   NAND2_X1 i_2959 (.A1(inputB[16]), .A2(inputA[12]), .ZN(n_3312));
   OAI21_X1 i_2960 (.A(n_3314), .B1(n_3462), .B2(n_3315), .ZN(n_3313));
   NAND2_X1 i_2961 (.A1(n_3462), .A2(n_3315), .ZN(n_3314));
   INV_X1 i_2962 (.A(n_3316), .ZN(n_3315));
   NAND2_X1 i_2963 (.A1(inputB[15]), .A2(inputA[13]), .ZN(n_3316));
   XOR2_X1 i_2964 (.A(n_3318), .B(n_3317), .Z(n_3038));
   NAND2_X1 i_2965 (.A1(inputB[13]), .A2(inputA[15]), .ZN(n_3317));
   NAND2_X1 i_2966 (.A1(n_3323), .A2(n_3319), .ZN(n_3318));
   NAND2_X1 i_2967 (.A1(n_3480), .A2(n_3322), .ZN(n_3319));
   AND2_X1 i_2968 (.A1(inputB[12]), .A2(inputA[17]), .ZN(n_3322));
   INV_X1 i_2969 (.A(n_3324), .ZN(n_3323));
   AOI22_X1 i_2970 (.A1(inputB[11]), .A2(inputA[17]), .B1(inputB[12]), .B2(
      inputA[16]), .ZN(n_3324));
   XOR2_X1 i_2971 (.A(n_3326), .B(n_3325), .Z(n_3052));
   NAND2_X1 i_2972 (.A1(inputB[7]), .A2(inputA[21]), .ZN(n_3325));
   OAI21_X1 i_2973 (.A(n_3329), .B1(n_3485), .B2(n_3330), .ZN(n_3326));
   NAND2_X1 i_2974 (.A1(n_3485), .A2(n_3330), .ZN(n_3329));
   INV_X1 i_2975 (.A(n_3331), .ZN(n_3330));
   NAND2_X1 i_2976 (.A1(inputB[6]), .A2(inputA[22]), .ZN(n_3331));
   XNOR2_X1 i_2977 (.A(n_3333), .B(n_3332), .ZN(n_3059));
   NAND2_X1 i_2978 (.A1(inputB[4]), .A2(inputA[24]), .ZN(n_3332));
   NOR2_X1 i_2979 (.A1(n_3335), .A2(n_3334), .ZN(n_3333));
   AOI21_X1 i_2980 (.A(n_3497), .B1(inputB[3]), .B2(inputA[25]), .ZN(n_3334));
   INV_X1 i_2981 (.A(n_3336), .ZN(n_3335));
   NAND3_X1 i_2982 (.A1(inputB[3]), .A2(inputA[25]), .A3(n_3497), .ZN(n_3336));
   AOI21_X1 i_2983 (.A(n_3337), .B1(n_3412), .B2(n_3411), .ZN(n_2919));
   NOR2_X1 i_2984 (.A1(n_3407), .A2(n_3403), .ZN(n_3337));
   INV_X1 i_2985 (.A(n_3338), .ZN(n_2928));
   AOI21_X1 i_2986 (.A(n_2925), .B1(n_2924), .B2(n_3371), .ZN(n_3338));
   OAI21_X1 i_2987 (.A(n_3360), .B1(n_3359), .B2(n_3356), .ZN(n_2856));
   OAI21_X1 i_2988 (.A(n_3432), .B1(n_3437), .B2(n_3427), .ZN(n_2863));
   OAI21_X1 i_2989 (.A(n_3385), .B1(n_3387), .B2(n_3382), .ZN(n_2877));
   OAI21_X1 i_2990 (.A(n_3458), .B1(n_3472), .B2(n_3453), .ZN(n_2884));
   OAI21_X1 i_2991 (.A(n_3380), .B1(n_3379), .B2(n_3376), .ZN(n_2898));
   OAI21_X1 i_2992 (.A(n_3484), .B1(n_3490), .B2(n_3482), .ZN(n_2905));
   XOR2_X1 i_2993 (.A(n_2994), .B(n_3339), .Z(n_2996));
   XOR2_X1 i_2994 (.A(n_2989), .B(n_3340), .Z(n_3339));
   XNOR2_X1 i_2995 (.A(n_2979), .B(n_3344), .ZN(n_3340));
   INV_X1 i_2996 (.A(n_3344), .ZN(n_3343));
   AOI21_X1 i_2997 (.A(n_2827), .B1(n_2826), .B2(n_3517), .ZN(n_3344));
   INV_X1 i_2998 (.A(n_3345), .ZN(n_2850));
   AOI21_X1 i_3000 (.A(n_2847), .B1(n_2846), .B2(n_3501), .ZN(n_3345));
   INV_X1 i_3001 (.A(n_3346), .ZN(n_2845));
   AOI21_X1 i_3002 (.A(n_2842), .B1(n_2841), .B2(n_3502), .ZN(n_3346));
   XNOR2_X1 i_3004 (.A(n_2984), .B(n_3350), .ZN(n_2986));
   INV_X1 i_3005 (.A(n_3350), .ZN(n_3347));
   AOI21_X1 i_3006 (.A(n_2832), .B1(n_2831), .B2(n_3503), .ZN(n_3350));
   INV_X1 i_3008 (.A(n_3351), .ZN(n_2840));
   AOI21_X1 i_3009 (.A(n_2837), .B1(n_2836), .B2(n_3512), .ZN(n_3351));
   XNOR2_X1 i_3010 (.A(n_2974), .B(n_3353), .ZN(n_2976));
   INV_X1 i_3012 (.A(n_3353), .ZN(n_3352));
   AOI21_X1 i_3013 (.A(n_2822), .B1(n_2821), .B2(n_3527), .ZN(n_3353));
   XOR2_X1 i_3014 (.A(n_2969), .B(n_3354), .Z(n_2971));
   XOR2_X1 i_3016 (.A(n_2949), .B(n_3355), .Z(n_3354));
   XOR2_X1 i_3017 (.A(n_3357), .B(n_3356), .Z(n_3355));
   NAND2_X1 i_3018 (.A1(inputB[27]), .A2(inputA[0]), .ZN(n_3356));
   NAND2_X1 i_3020 (.A1(n_3360), .A2(n_3358), .ZN(n_3357));
   INV_X1 i_3021 (.A(n_3359), .ZN(n_3358));
   AOI22_X1 i_3022 (.A1(inputB[25]), .A2(inputA[2]), .B1(inputB[26]), .B2(
      inputA[1]), .ZN(n_3359));
   NAND2_X1 i_3024 (.A1(n_3597), .A2(n_3361), .ZN(n_3360));
   INV_X1 i_3025 (.A(n_3364), .ZN(n_3361));
   NAND2_X1 i_3026 (.A1(inputB[26]), .A2(inputA[2]), .ZN(n_3364));
   XOR2_X1 i_3028 (.A(n_2964), .B(n_3365), .Z(n_2966));
   XNOR2_X1 i_3029 (.A(n_2934), .B(n_3367), .ZN(n_3365));
   INV_X1 i_3030 (.A(n_3367), .ZN(n_3366));
   AOI21_X1 i_3032 (.A(n_2777), .B1(n_2776), .B2(n_3505), .ZN(n_3367));
   XOR2_X1 i_3033 (.A(n_2954), .B(n_3368), .Z(n_2956));
   XOR2_X1 i_3034 (.A(n_2924), .B(n_3371), .Z(n_3368));
   NAND2_X1 i_3036 (.A1(n_3644), .A2(n_3372), .ZN(n_3371));
   NAND2_X1 i_3037 (.A1(n_3643), .A2(n_3638), .ZN(n_3372));
   XNOR2_X1 i_3038 (.A(n_2959), .B(n_3374), .ZN(n_2961));
   INV_X1 i_3040 (.A(n_3374), .ZN(n_3373));
   AOI21_X1 i_3041 (.A(n_2797), .B1(n_2796), .B2(n_3518), .ZN(n_3374));
   XOR2_X1 i_3042 (.A(n_2939), .B(n_3375), .Z(n_2941));
   XOR2_X1 i_3044 (.A(n_3377), .B(n_3376), .Z(n_3375));
   NAND2_X1 i_3045 (.A1(inputB[9]), .A2(inputA[18]), .ZN(n_3376));
   NAND2_X1 i_3046 (.A1(n_3380), .A2(n_3378), .ZN(n_3377));
   INV_X1 i_3048 (.A(n_3379), .ZN(n_3378));
   AOI22_X1 i_3049 (.A1(inputB[7]), .A2(inputA[20]), .B1(inputB[8]), .B2(
      inputA[19]), .ZN(n_3379));
   NAND3_X1 i_3050 (.A1(inputB[8]), .A2(inputA[20]), .A3(n_3655), .ZN(n_3380));
   XOR2_X1 i_3052 (.A(n_2944), .B(n_3381), .Z(n_2946));
   XOR2_X1 i_3053 (.A(n_3384), .B(n_3382), .Z(n_3381));
   NAND2_X1 i_3054 (.A1(inputB[18]), .A2(inputA[9]), .ZN(n_3382));
   NAND2_X1 i_3056 (.A1(n_3386), .A2(n_3385), .ZN(n_3384));
   NAND3_X1 i_3057 (.A1(inputB[17]), .A2(inputA[11]), .A3(n_3637), .ZN(n_3385));
   INV_X1 i_3058 (.A(n_3387), .ZN(n_3386));
   AOI22_X1 i_3060 (.A1(inputB[16]), .A2(inputA[11]), .B1(inputB[17]), .B2(
      inputA[10]), .ZN(n_3387));
   INV_X1 i_3061 (.A(n_3388), .ZN(n_2815));
   AOI21_X1 i_3062 (.A(n_2812), .B1(n_2811), .B2(n_3504), .ZN(n_3388));
   INV_X1 i_3064 (.A(n_3392), .ZN(n_2820));
   AOI21_X1 i_3065 (.A(n_2817), .B1(n_2816), .B2(n_3533), .ZN(n_3392));
   INV_X1 i_3066 (.A(n_3396), .ZN(n_2810));
   AOI21_X1 i_3068 (.A(n_2807), .B1(n_2806), .B2(n_3546), .ZN(n_3396));
   INV_X1 i_3069 (.A(n_3397), .ZN(n_2795));
   AOI21_X1 i_3070 (.A(n_2792), .B1(n_2791), .B2(n_3551), .ZN(n_3397));
   INV_X1 i_3071 (.A(n_3402), .ZN(n_2805));
   AOI21_X1 i_3072 (.A(n_2802), .B1(n_2801), .B2(n_3537), .ZN(n_3402));
   XOR2_X1 i_3073 (.A(n_3406), .B(n_3403), .Z(n_2918));
   AND2_X1 i_3074 (.A1(inputB[0]), .A2(inputA[27]), .ZN(n_3403));
   AOI21_X1 i_3075 (.A(n_3407), .B1(n_3412), .B2(n_3411), .ZN(n_3406));
   NOR2_X1 i_3076 (.A1(n_3412), .A2(n_3411), .ZN(n_3407));
   AOI22_X1 i_3077 (.A1(n_3679), .A2(n_3662), .B1(n_3659), .B2(n_3657), .ZN(
      n_3411));
   INV_X1 i_3078 (.A(n_3413), .ZN(n_3412));
   OAI21_X1 i_3079 (.A(n_3554), .B1(n_3558), .B2(n_3552), .ZN(n_3413));
   XOR2_X1 i_3080 (.A(n_2929), .B(n_3417), .Z(n_2931));
   OAI21_X1 i_3081 (.A(n_3608), .B1(n_3618), .B2(n_3598), .ZN(n_3417));
   INV_X1 i_3082 (.A(n_3422), .ZN(n_2790));
   AOI21_X1 i_3083 (.A(n_2787), .B1(n_2786), .B2(n_3573), .ZN(n_3422));
   XOR2_X1 i_3084 (.A(n_3431), .B(n_3427), .Z(n_2862));
   NAND2_X1 i_3085 (.A1(inputB[24]), .A2(inputA[3]), .ZN(n_3427));
   NAND2_X1 i_3086 (.A1(n_3433), .A2(n_3432), .ZN(n_3431));
   NAND4_X1 i_3087 (.A1(inputB[22]), .A2(inputA[5]), .A3(inputB[23]), .A4(
      inputA[4]), .ZN(n_3432));
   INV_X1 i_3088 (.A(n_3437), .ZN(n_3433));
   AOI22_X1 i_3089 (.A1(inputB[22]), .A2(inputA[5]), .B1(inputB[23]), .B2(
      inputA[4]), .ZN(n_3437));
   XOR2_X1 i_3090 (.A(n_3442), .B(n_3441), .Z(n_2869));
   NAND2_X1 i_3091 (.A1(inputB[21]), .A2(inputA[6]), .ZN(n_3441));
   OAI21_X1 i_3092 (.A(n_3443), .B1(n_3544), .B2(n_3447), .ZN(n_3442));
   NAND2_X1 i_3093 (.A1(n_3544), .A2(n_3447), .ZN(n_3443));
   INV_X1 i_3094 (.A(n_3452), .ZN(n_3447));
   NAND2_X1 i_3095 (.A1(inputB[20]), .A2(inputA[7]), .ZN(n_3452));
   XOR2_X1 i_3096 (.A(n_3457), .B(n_3453), .Z(n_2883));
   NAND2_X1 i_3097 (.A1(inputB[15]), .A2(inputA[12]), .ZN(n_3453));
   NAND2_X1 i_3098 (.A1(n_3467), .A2(n_3458), .ZN(n_3457));
   NAND2_X1 i_3099 (.A1(n_3647), .A2(n_3462), .ZN(n_3458));
   INV_X1 i_3100 (.A(n_3466), .ZN(n_3462));
   NAND2_X1 i_3101 (.A1(inputB[14]), .A2(inputA[14]), .ZN(n_3466));
   INV_X1 i_3102 (.A(n_3472), .ZN(n_3467));
   AOI22_X1 i_3103 (.A1(inputB[13]), .A2(inputA[14]), .B1(inputB[14]), .B2(
      inputA[13]), .ZN(n_3472));
   XOR2_X1 i_3104 (.A(n_3478), .B(n_3476), .Z(n_2890));
   NAND2_X1 i_3105 (.A1(inputB[12]), .A2(inputA[15]), .ZN(n_3476));
   OAI21_X1 i_3106 (.A(n_3479), .B1(n_3525), .B2(n_3480), .ZN(n_3478));
   NAND2_X1 i_3107 (.A1(n_3525), .A2(n_3480), .ZN(n_3479));
   INV_X1 i_3108 (.A(n_3481), .ZN(n_3480));
   NAND2_X1 i_3109 (.A1(inputB[11]), .A2(inputA[16]), .ZN(n_3481));
   XOR2_X1 i_3110 (.A(n_3483), .B(n_3482), .Z(n_2904));
   NAND2_X1 i_3111 (.A1(inputB[6]), .A2(inputA[21]), .ZN(n_3482));
   NAND2_X1 i_3112 (.A1(n_3489), .A2(n_3484), .ZN(n_3483));
   NAND2_X1 i_3113 (.A1(n_3662), .A2(n_3485), .ZN(n_3484));
   INV_X1 i_3114 (.A(n_3488), .ZN(n_3485));
   NAND2_X1 i_3115 (.A1(inputB[5]), .A2(inputA[23]), .ZN(n_3488));
   INV_X1 i_3116 (.A(n_3490), .ZN(n_3489));
   AOI22_X1 i_3117 (.A1(inputB[4]), .A2(inputA[23]), .B1(inputB[5]), .B2(
      inputA[22]), .ZN(n_3490));
   XOR2_X1 i_3118 (.A(n_3492), .B(n_3491), .Z(n_2911));
   NAND2_X1 i_3119 (.A1(inputB[3]), .A2(inputA[24]), .ZN(n_3491));
   NAND2_X1 i_3120 (.A1(n_3496), .A2(n_3493), .ZN(n_3492));
   INV_X1 i_3121 (.A(n_3495), .ZN(n_3493));
   AOI22_X1 i_3122 (.A1(inputB[1]), .A2(inputA[26]), .B1(inputB[2]), .B2(
      inputA[25]), .ZN(n_3495));
   NAND3_X1 i_3123 (.A1(inputB[1]), .A2(inputA[25]), .A3(n_3497), .ZN(n_3496));
   AND2_X1 i_3124 (.A1(inputB[2]), .A2(inputA[26]), .ZN(n_3497));
   INV_X1 i_3125 (.A(n_3498), .ZN(n_2785));
   AOI21_X1 i_3126 (.A(n_2782), .B1(n_2781), .B2(n_3568), .ZN(n_3498));
   OAI21_X1 i_3127 (.A(n_3587), .B1(n_3593), .B2(n_3583), .ZN(n_2716));
   OAI21_X1 i_3128 (.A(n_3543), .B1(n_3541), .B2(n_3538), .ZN(n_2730));
   OAI21_X1 i_3129 (.A(n_3627), .B1(n_3633), .B2(n_3619), .ZN(n_2737));
   OAI21_X1 i_3130 (.A(n_3524), .B1(n_3523), .B2(n_3519), .ZN(n_2751));
   NAND2_X1 i_3131 (.A1(n_3654), .A2(n_3499), .ZN(n_2758));
   NAND2_X1 i_3132 (.A1(n_3652), .A2(n_3650), .ZN(n_3499));
   XOR2_X1 i_3133 (.A(n_2846), .B(n_3501), .Z(n_2848));
   XOR2_X1 i_3134 (.A(n_2841), .B(n_3502), .Z(n_3501));
   XOR2_X1 i_3135 (.A(n_2831), .B(n_3503), .Z(n_3502));
   XOR2_X1 i_3136 (.A(n_2811), .B(n_3504), .Z(n_3503));
   XOR2_X1 i_3137 (.A(n_2776), .B(n_3505), .Z(n_3504));
   AOI22_X1 i_3138 (.A1(n_3902), .A2(n_3766), .B1(n_3764), .B2(n_3759), .ZN(
      n_3505));
   INV_X1 i_3139 (.A(n_3506), .ZN(n_2710));
   AOI21_X1 i_3140 (.A(n_2707), .B1(n_2706), .B2(n_3509), .ZN(n_3506));
   XOR2_X1 i_3141 (.A(n_2701), .B(n_3511), .Z(n_3509));
   INV_X1 i_3142 (.A(n_3510), .ZN(n_2705));
   AOI21_X1 i_3143 (.A(n_2702), .B1(n_2701), .B2(n_3511), .ZN(n_3510));
   XOR2_X1 i_3144 (.A(n_2691), .B(n_3514), .Z(n_3511));
   XNOR2_X1 i_3145 (.A(n_2836), .B(n_3513), .ZN(n_2838));
   INV_X1 i_3147 (.A(n_3513), .ZN(n_3512));
   AOI21_X1 i_3148 (.A(n_2692), .B1(n_2691), .B2(n_3514), .ZN(n_3513));
   XOR2_X1 i_3149 (.A(n_2671), .B(n_3531), .Z(n_3514));
   INV_X1 i_3151 (.A(n_3516), .ZN(n_2700));
   AOI21_X1 i_3152 (.A(n_2697), .B1(n_2696), .B2(n_3667), .ZN(n_3516));
   XOR2_X1 i_3153 (.A(n_2826), .B(n_3517), .Z(n_2828));
   XOR2_X1 i_3155 (.A(n_2796), .B(n_3518), .Z(n_3517));
   XOR2_X1 i_3156 (.A(n_3520), .B(n_3519), .Z(n_3518));
   NAND2_X1 i_3157 (.A1(inputB[11]), .A2(inputA[15]), .ZN(n_3519));
   NAND2_X1 i_3159 (.A1(n_3524), .A2(n_3522), .ZN(n_3520));
   INV_X1 i_3160 (.A(n_3523), .ZN(n_3522));
   AOI22_X1 i_3161 (.A1(inputB[9]), .A2(inputA[17]), .B1(inputB[10]), .B2(
      inputA[16]), .ZN(n_3523));
   NAND2_X1 i_3163 (.A1(n_3765), .A2(n_3525), .ZN(n_3524));
   INV_X1 i_3164 (.A(n_3526), .ZN(n_3525));
   NAND2_X1 i_3165 (.A1(inputB[10]), .A2(inputA[17]), .ZN(n_3526));
   XNOR2_X1 i_3167 (.A(n_2821), .B(n_3530), .ZN(n_2823));
   INV_X1 i_3168 (.A(n_3530), .ZN(n_3527));
   AOI21_X1 i_3169 (.A(n_2672), .B1(n_2671), .B2(n_3531), .ZN(n_3530));
   XOR2_X1 i_3171 (.A(n_2641), .B(n_3665), .Z(n_3531));
   INV_X1 i_3172 (.A(n_3532), .ZN(n_2690));
   AOI21_X1 i_3173 (.A(n_2687), .B1(n_2686), .B2(n_3671), .ZN(n_3532));
   XNOR2_X1 i_3175 (.A(n_2816), .B(n_3534), .ZN(n_2818));
   INV_X1 i_3176 (.A(n_3534), .ZN(n_3533));
   AOI21_X1 i_3177 (.A(n_2657), .B1(n_2656), .B2(n_3672), .ZN(n_3534));
   INV_X1 i_3179 (.A(n_3535), .ZN(n_2685));
   AOI21_X1 i_3180 (.A(n_2682), .B1(n_2681), .B2(n_3684), .ZN(n_3535));
   XOR2_X1 i_3181 (.A(n_2801), .B(n_3537), .Z(n_2803));
   XOR2_X1 i_3183 (.A(n_3539), .B(n_3538), .Z(n_3537));
   NAND2_X1 i_3184 (.A1(inputB[20]), .A2(inputA[6]), .ZN(n_3538));
   NAND2_X1 i_3185 (.A1(n_3543), .A2(n_3540), .ZN(n_3539));
   INV_X1 i_3187 (.A(n_3541), .ZN(n_3540));
   AOI22_X1 i_3188 (.A1(inputB[18]), .A2(inputA[8]), .B1(inputB[19]), .B2(
      inputA[7]), .ZN(n_3541));
   NAND2_X1 i_3189 (.A1(n_3740), .A2(n_3544), .ZN(n_3543));
   INV_X1 i_3191 (.A(n_3545), .ZN(n_3544));
   NAND2_X1 i_3192 (.A1(inputB[19]), .A2(inputA[8]), .ZN(n_3545));
   XNOR2_X1 i_3193 (.A(n_2806), .B(n_3547), .ZN(n_2808));
   INV_X1 i_3195 (.A(n_3547), .ZN(n_3546));
   AOI21_X1 i_3196 (.A(n_2652), .B1(n_2651), .B2(n_3711), .ZN(n_3547));
   INV_X1 i_3197 (.A(n_3548), .ZN(n_2680));
   AOI21_X1 i_3199 (.A(n_2677), .B1(n_2676), .B2(n_3687), .ZN(n_3548));
   XOR2_X1 i_3200 (.A(n_2791), .B(n_3551), .Z(n_2793));
   XOR2_X1 i_3201 (.A(n_3553), .B(n_3552), .Z(n_3551));
   NAND2_X1 i_3203 (.A1(inputB[2]), .A2(inputA[24]), .ZN(n_3552));
   NAND2_X1 i_3204 (.A1(n_3557), .A2(n_3554), .ZN(n_3553));
   NAND3_X1 i_3205 (.A1(inputB[1]), .A2(inputA[26]), .A3(n_3806), .ZN(n_3554));
   INV_X1 i_3207 (.A(n_3558), .ZN(n_3557));
   AOI22_X1 i_3208 (.A1(inputB[0]), .A2(inputA[26]), .B1(inputB[1]), .B2(
      inputA[25]), .ZN(n_3558));
   INV_X1 i_3209 (.A(n_3559), .ZN(n_2665));
   AOI21_X1 i_3211 (.A(n_2662), .B1(n_2661), .B2(n_3691), .ZN(n_3559));
   INV_X1 i_3212 (.A(n_3563), .ZN(n_2670));
   AOI21_X1 i_3213 (.A(n_2667), .B1(n_2666), .B2(n_3700), .ZN(n_3563));
   XOR2_X1 i_3215 (.A(n_2781), .B(n_3568), .Z(n_2783));
   OAI21_X1 i_3216 (.A(n_3731), .B1(n_3739), .B2(n_3729), .ZN(n_3568));
   XNOR2_X1 i_3217 (.A(n_2786), .B(n_3578), .ZN(n_2788));
   INV_X1 i_3218 (.A(n_3578), .ZN(n_3573));
   AOI21_X1 i_3219 (.A(n_2647), .B1(n_2646), .B2(n_3715), .ZN(n_3578));
   XOR2_X1 i_3220 (.A(n_3584), .B(n_3583), .Z(n_2715));
   NAND2_X1 i_3221 (.A1(inputB[26]), .A2(inputA[0]), .ZN(n_3583));
   NAND2_X1 i_3222 (.A1(n_3588), .A2(n_3587), .ZN(n_3584));
   NAND3_X1 i_3223 (.A1(inputB[24]), .A2(inputA[2]), .A3(n_3597), .ZN(n_3587));
   INV_X1 i_3224 (.A(n_3593), .ZN(n_3588));
   AOI21_X1 i_3225 (.A(n_3597), .B1(inputB[24]), .B2(inputA[2]), .ZN(n_3593));
   AND2_X1 i_3226 (.A1(inputB[25]), .A2(inputA[1]), .ZN(n_3597));
   XOR2_X1 i_3227 (.A(n_3603), .B(n_3598), .Z(n_2722));
   NAND2_X1 i_3228 (.A1(inputB[23]), .A2(inputA[3]), .ZN(n_3598));
   NAND2_X1 i_3229 (.A1(n_3613), .A2(n_3608), .ZN(n_3603));
   NAND3_X1 i_3230 (.A1(inputB[22]), .A2(inputA[4]), .A3(n_3706), .ZN(n_3608));
   INV_X1 i_3231 (.A(n_3618), .ZN(n_3613));
   AOI21_X1 i_3232 (.A(n_3706), .B1(inputB[22]), .B2(inputA[4]), .ZN(n_3618));
   XOR2_X1 i_3233 (.A(n_3623), .B(n_3619), .Z(n_2736));
   NAND2_X1 i_3234 (.A1(inputB[17]), .A2(inputA[9]), .ZN(n_3619));
   NAND2_X1 i_3235 (.A1(n_3628), .A2(n_3627), .ZN(n_3623));
   NAND3_X1 i_3236 (.A1(inputB[15]), .A2(inputA[11]), .A3(n_3637), .ZN(n_3627));
   INV_X1 i_3237 (.A(n_3633), .ZN(n_3628));
   AOI21_X1 i_3238 (.A(n_3637), .B1(inputB[15]), .B2(inputA[11]), .ZN(n_3633));
   AND2_X1 i_3239 (.A1(inputB[16]), .A2(inputA[10]), .ZN(n_3637));
   XOR2_X1 i_3240 (.A(n_3639), .B(n_3638), .Z(n_2743));
   AND2_X1 i_3241 (.A1(inputB[14]), .A2(inputA[12]), .ZN(n_3638));
   AND2_X1 i_3242 (.A1(n_3644), .A2(n_3643), .ZN(n_3639));
   NAND2_X1 i_3243 (.A1(n_3699), .A2(n_3648), .ZN(n_3643));
   NAND2_X1 i_3244 (.A1(n_3698), .A2(n_3647), .ZN(n_3644));
   INV_X1 i_3245 (.A(n_3648), .ZN(n_3647));
   NAND2_X1 i_3246 (.A1(inputB[13]), .A2(inputA[13]), .ZN(n_3648));
   XOR2_X1 i_3247 (.A(n_3651), .B(n_3650), .Z(n_2757));
   AND2_X1 i_3248 (.A1(inputB[8]), .A2(inputA[18]), .ZN(n_3650));
   AND2_X1 i_3249 (.A1(n_3654), .A2(n_3652), .ZN(n_3651));
   NAND2_X1 i_3250 (.A1(n_3784), .A2(n_3656), .ZN(n_3652));
   NAND2_X1 i_3251 (.A1(n_3781), .A2(n_3655), .ZN(n_3654));
   INV_X1 i_3252 (.A(n_3656), .ZN(n_3655));
   NAND2_X1 i_3253 (.A1(inputB[7]), .A2(inputA[19]), .ZN(n_3656));
   XOR2_X1 i_3254 (.A(n_3658), .B(n_3657), .Z(n_2764));
   AND2_X1 i_3255 (.A1(inputB[5]), .A2(inputA[21]), .ZN(n_3657));
   AOI22_X1 i_3256 (.A1(n_3679), .A2(n_3662), .B1(n_3680), .B2(n_3663), .ZN(
      n_3658));
   NAND2_X1 i_3257 (.A1(n_3680), .A2(n_3663), .ZN(n_3659));
   INV_X1 i_3258 (.A(n_3663), .ZN(n_3662));
   NAND2_X1 i_3259 (.A1(inputB[4]), .A2(inputA[22]), .ZN(n_3663));
   OAI21_X1 i_3260 (.A(n_3796), .B1(n_3800), .B2(n_3794), .ZN(n_2635));
   INV_X1 i_3261 (.A(n_3664), .ZN(n_2645));
   AOI21_X1 i_3262 (.A(n_2642), .B1(n_2641), .B2(n_3665), .ZN(n_3664));
   AOI21_X1 i_3263 (.A(n_3841), .B1(n_3840), .B2(n_3837), .ZN(n_3665));
   OAI21_X1 i_3264 (.A(n_3720), .B1(n_3725), .B2(n_3718), .ZN(n_2580));
   OAI21_X1 i_3265 (.A(n_3705), .B1(n_3708), .B2(n_3701), .ZN(n_2587));
   OAI21_X1 i_3266 (.A(n_3750), .B1(n_3756), .B2(n_3744), .ZN(n_2601));
   OAI21_X1 i_3267 (.A(n_3697), .B1(n_3696), .B2(n_3692), .ZN(n_2608));
   OAI21_X1 i_3268 (.A(n_3780), .B1(n_3790), .B2(n_3770), .ZN(n_2622));
   OAI21_X1 i_3269 (.A(n_3678), .B1(n_3677), .B2(n_3673), .ZN(n_2629));
   INV_X1 i_3270 (.A(n_3666), .ZN(n_2574));
   AOI21_X1 i_3271 (.A(n_2571), .B1(n_2570), .B2(n_3817), .ZN(n_3666));
   XNOR2_X1 i_3272 (.A(n_2696), .B(n_3669), .ZN(n_2698));
   INV_X1 i_3273 (.A(n_3669), .ZN(n_3667));
   AOI21_X1 i_3274 (.A(n_2556), .B1(n_2555), .B2(n_3819), .ZN(n_3669));
   INV_X1 i_3275 (.A(n_3670), .ZN(n_2569));
   AOI21_X1 i_3276 (.A(n_2566), .B1(n_2565), .B2(n_3818), .ZN(n_3670));
   XOR2_X1 i_3277 (.A(n_2686), .B(n_3671), .Z(n_2688));
   XOR2_X1 i_3278 (.A(n_2656), .B(n_3672), .Z(n_3671));
   XOR2_X1 i_3279 (.A(n_3675), .B(n_3673), .Z(n_3672));
   NAND2_X1 i_3280 (.A1(inputB[4]), .A2(inputA[21]), .ZN(n_3673));
   NAND2_X1 i_3281 (.A1(n_3678), .A2(n_3676), .ZN(n_3675));
   INV_X1 i_3282 (.A(n_3677), .ZN(n_3676));
   AOI22_X1 i_3283 (.A1(inputB[2]), .A2(inputA[23]), .B1(inputB[3]), .B2(
      inputA[22]), .ZN(n_3677));
   NAND3_X1 i_3284 (.A1(inputB[2]), .A2(inputA[22]), .A3(n_3679), .ZN(n_3678));
   INV_X1 i_3285 (.A(n_3680), .ZN(n_3679));
   NAND2_X1 i_3286 (.A1(inputB[3]), .A2(inputA[23]), .ZN(n_3680));
   INV_X1 i_3287 (.A(n_3683), .ZN(n_2564));
   AOI21_X1 i_3288 (.A(n_2561), .B1(n_2560), .B2(n_3831), .ZN(n_3683));
   XNOR2_X1 i_3289 (.A(n_2681), .B(n_3685), .ZN(n_2683));
   INV_X1 i_3290 (.A(n_3685), .ZN(n_3684));
   AOI21_X1 i_3291 (.A(n_2536), .B1(n_2535), .B2(n_3847), .ZN(n_3685));
   INV_X1 i_3292 (.A(n_3686), .ZN(n_2554));
   AOI21_X1 i_3293 (.A(n_2551), .B1(n_2550), .B2(n_3833), .ZN(n_3686));
   XNOR2_X1 i_3295 (.A(n_2676), .B(n_3688), .ZN(n_2678));
   INV_X1 i_3296 (.A(n_3688), .ZN(n_3687));
   AOI21_X1 i_3297 (.A(n_2521), .B1(n_2520), .B2(n_3821), .ZN(n_3688));
   INV_X1 i_3299 (.A(n_3690), .ZN(n_2549));
   AOI21_X1 i_3300 (.A(n_2546), .B1(n_2545), .B2(n_3820), .ZN(n_3690));
   XOR2_X1 i_3301 (.A(n_2661), .B(n_3691), .Z(n_2663));
   XOR2_X1 i_3303 (.A(n_3693), .B(n_3692), .Z(n_3691));
   NAND2_X1 i_3304 (.A1(inputB[13]), .A2(inputA[12]), .ZN(n_3692));
   NAND2_X1 i_3305 (.A1(n_3697), .A2(n_3694), .ZN(n_3693));
   INV_X1 i_3307 (.A(n_3696), .ZN(n_3694));
   AOI22_X1 i_3308 (.A1(inputB[11]), .A2(inputA[14]), .B1(inputB[12]), .B2(
      inputA[13]), .ZN(n_3696));
   NAND3_X1 i_3309 (.A1(inputB[11]), .A2(inputA[13]), .A3(n_3698), .ZN(n_3697));
   INV_X1 i_3311 (.A(n_3699), .ZN(n_3698));
   NAND2_X1 i_3312 (.A1(inputB[12]), .A2(inputA[14]), .ZN(n_3699));
   XOR2_X1 i_3313 (.A(n_2666), .B(n_3700), .Z(n_2668));
   XOR2_X1 i_3315 (.A(n_3704), .B(n_3701), .Z(n_3700));
   NAND2_X1 i_3316 (.A1(inputB[22]), .A2(inputA[3]), .ZN(n_3701));
   NAND2_X1 i_3317 (.A1(n_3707), .A2(n_3705), .ZN(n_3704));
   NAND3_X1 i_3319 (.A1(inputB[20]), .A2(inputA[4]), .A3(n_3706), .ZN(n_3705));
   AND2_X1 i_3320 (.A1(inputB[21]), .A2(inputA[5]), .ZN(n_3706));
   INV_X1 i_3321 (.A(n_3708), .ZN(n_3707));
   AOI22_X1 i_3323 (.A1(inputB[20]), .A2(inputA[5]), .B1(inputB[21]), .B2(
      inputA[4]), .ZN(n_3708));
   INV_X1 i_3324 (.A(n_3709), .ZN(n_2544));
   AOI21_X1 i_3325 (.A(n_2541), .B1(n_2540), .B2(n_3844), .ZN(n_3709));
   XNOR2_X1 i_3327 (.A(n_2651), .B(n_3712), .ZN(n_2653));
   INV_X1 i_3328 (.A(n_3712), .ZN(n_3711));
   AOI21_X1 i_3329 (.A(n_2511), .B1(n_2510), .B2(n_3868), .ZN(n_3712));
   INV_X1 i_3331 (.A(n_3713), .ZN(n_2529));
   AOI21_X1 i_3332 (.A(n_2526), .B1(n_2525), .B2(n_3836), .ZN(n_3713));
   INV_X1 i_3333 (.A(n_3714), .ZN(n_2534));
   AOI21_X1 i_3335 (.A(n_2531), .B1(n_2530), .B2(n_3851), .ZN(n_3714));
   XOR2_X1 i_3336 (.A(n_2646), .B(n_3715), .Z(n_2648));
   OAI21_X1 i_3337 (.A(n_3854), .B1(n_3858), .B2(n_3852), .ZN(n_3715));
   XOR2_X1 i_3339 (.A(n_3719), .B(n_3718), .Z(n_2579));
   NAND2_X1 i_3340 (.A1(inputB[25]), .A2(inputA[0]), .ZN(n_3718));
   NAND2_X1 i_3341 (.A1(n_3721), .A2(n_3720), .ZN(n_3719));
   NAND4_X1 i_3343 (.A1(inputB[23]), .A2(inputA[2]), .A3(inputB[24]), .A4(
      inputA[1]), .ZN(n_3720));
   INV_X1 i_3344 (.A(n_3725), .ZN(n_3721));
   AOI22_X1 i_3345 (.A1(inputB[23]), .A2(inputA[2]), .B1(inputB[24]), .B2(
      inputA[1]), .ZN(n_3725));
   XOR2_X1 i_3347 (.A(n_3730), .B(n_3729), .Z(n_2593));
   NAND2_X1 i_3348 (.A1(inputB[19]), .A2(inputA[6]), .ZN(n_3729));
   NAND2_X1 i_3349 (.A1(n_3735), .A2(n_3731), .ZN(n_3730));
   NAND3_X1 i_3351 (.A1(inputB[17]), .A2(inputA[8]), .A3(n_3740), .ZN(n_3731));
   INV_X1 i_3352 (.A(n_3739), .ZN(n_3735));
   AOI21_X1 i_3353 (.A(n_3740), .B1(inputB[17]), .B2(inputA[8]), .ZN(n_3739));
   AND2_X1 i_3355 (.A1(inputB[18]), .A2(inputA[7]), .ZN(n_3740));
   XOR2_X1 i_3356 (.A(n_3745), .B(n_3744), .Z(n_2600));
   NAND2_X1 i_3357 (.A1(inputB[16]), .A2(inputA[9]), .ZN(n_3744));
   NAND2_X1 i_3359 (.A1(n_3755), .A2(n_3750), .ZN(n_3745));
   NAND4_X1 i_3360 (.A1(inputB[14]), .A2(inputA[11]), .A3(inputB[15]), .A4(
      inputA[10]), .ZN(n_3750));
   INV_X1 i_3361 (.A(n_3756), .ZN(n_3755));
   AOI22_X1 i_3363 (.A1(inputB[14]), .A2(inputA[11]), .B1(inputB[15]), .B2(
      inputA[10]), .ZN(n_3756));
   XOR2_X1 i_3364 (.A(n_3760), .B(n_3759), .Z(n_2614));
   NAND2_X1 i_3365 (.A1(inputB[10]), .A2(inputA[15]), .ZN(n_3759));
   OAI21_X1 i_3367 (.A(n_3764), .B1(n_3897), .B2(n_3765), .ZN(n_3760));
   NAND2_X1 i_3368 (.A1(n_3897), .A2(n_3765), .ZN(n_3764));
   INV_X1 i_3369 (.A(n_3766), .ZN(n_3765));
   NAND2_X1 i_3370 (.A1(inputB[9]), .A2(inputA[16]), .ZN(n_3766));
   XOR2_X1 i_3371 (.A(n_3775), .B(n_3770), .Z(n_2621));
   NAND2_X1 i_3372 (.A1(inputB[7]), .A2(inputA[18]), .ZN(n_3770));
   NAND2_X1 i_3373 (.A1(n_3785), .A2(n_3780), .ZN(n_3775));
   NAND2_X1 i_3374 (.A1(n_3917), .A2(n_3781), .ZN(n_3780));
   INV_X1 i_3375 (.A(n_3784), .ZN(n_3781));
   NAND2_X1 i_3376 (.A1(inputB[6]), .A2(inputA[20]), .ZN(n_3784));
   INV_X1 i_3377 (.A(n_3790), .ZN(n_3785));
   AOI22_X1 i_3378 (.A1(inputB[5]), .A2(inputA[20]), .B1(inputB[6]), .B2(
      inputA[19]), .ZN(n_3790));
   XOR2_X1 i_3379 (.A(n_3795), .B(n_3794), .Z(n_2634));
   NAND2_X1 i_3380 (.A1(inputB[1]), .A2(inputA[24]), .ZN(n_3794));
   OAI21_X1 i_3381 (.A(n_3796), .B1(n_3806), .B2(n_3805), .ZN(n_3795));
   NAND2_X1 i_3382 (.A1(n_3806), .A2(n_3805), .ZN(n_3796));
   NOR2_X1 i_3383 (.A1(n_3806), .A2(n_3805), .ZN(n_3800));
   OAI21_X1 i_3384 (.A(n_3826), .B1(n_3825), .B2(n_3822), .ZN(n_3805));
   AND2_X1 i_3385 (.A1(inputB[0]), .A2(inputA[25]), .ZN(n_3806));
   AOI21_X1 i_3386 (.A(n_3810), .B1(n_3866), .B2(n_3865), .ZN(n_2505));
   NOR2_X1 i_3387 (.A1(n_3864), .A2(n_3862), .ZN(n_3810));
   INV_X1 i_3388 (.A(n_3815), .ZN(n_2519));
   AOI21_X1 i_3389 (.A(n_2516), .B1(n_2515), .B2(n_3850), .ZN(n_3815));
   OAI21_X1 i_3390 (.A(n_3874), .B1(n_3878), .B2(n_3872), .ZN(n_2449));
   OAI21_X1 i_3391 (.A(n_3881), .B1(n_3883), .B2(n_3879), .ZN(n_2463));
   OAI21_X1 i_3392 (.A(n_3886), .B1(n_3888), .B2(n_3884), .ZN(n_2470));
   OAI21_X1 i_3393 (.A(n_3896), .B1(n_3911), .B2(n_3892), .ZN(n_2484));
   AOI22_X1 i_3394 (.A1(n_3995), .A2(n_3922), .B1(n_3916), .B2(n_3912), .ZN(
      n_2491));
   XOR2_X1 i_3395 (.A(n_2570), .B(n_3817), .Z(n_2572));
   XOR2_X1 i_3396 (.A(n_2565), .B(n_3818), .Z(n_3817));
   XOR2_X1 i_3397 (.A(n_2555), .B(n_3819), .Z(n_3818));
   XOR2_X1 i_3398 (.A(n_2545), .B(n_3820), .Z(n_3819));
   XOR2_X1 i_3399 (.A(n_2520), .B(n_3821), .Z(n_3820));
   XOR2_X1 i_3400 (.A(n_3823), .B(n_3822), .Z(n_3821));
   NAND2_X1 i_3401 (.A1(inputB[3]), .A2(inputA[21]), .ZN(n_3822));
   NAND2_X1 i_3402 (.A1(n_3826), .A2(n_3824), .ZN(n_3823));
   INV_X1 i_3403 (.A(n_3825), .ZN(n_3824));
   AOI22_X1 i_3404 (.A1(inputB[1]), .A2(inputA[23]), .B1(inputB[2]), .B2(
      inputA[22]), .ZN(n_3825));
   NAND3_X1 i_3405 (.A1(inputB[2]), .A2(inputA[23]), .A3(n_4146), .ZN(n_3826));
   INV_X1 i_3406 (.A(n_3829), .ZN(n_2443));
   AOI21_X1 i_3407 (.A(n_2440), .B1(n_2439), .B2(n_3933), .ZN(n_3829));
   INV_X1 i_3408 (.A(n_3830), .ZN(n_2438));
   AOI21_X1 i_3409 (.A(n_2435), .B1(n_2434), .B2(n_3936), .ZN(n_3830));
   XNOR2_X1 i_3410 (.A(n_2560), .B(n_3832), .ZN(n_2562));
   INV_X1 i_3411 (.A(n_3832), .ZN(n_3831));
   AOI21_X1 i_3412 (.A(n_2425), .B1(n_2424), .B2(n_3937), .ZN(n_3832));
   XOR2_X1 i_3413 (.A(n_2550), .B(n_3833), .Z(n_2552));
   XOR2_X1 i_3414 (.A(n_2525), .B(n_3836), .Z(n_3833));
   XNOR2_X1 i_3415 (.A(n_3838), .B(n_3837), .ZN(n_3836));
   NAND2_X1 i_3416 (.A1(inputB[12]), .A2(inputA[12]), .ZN(n_3837));
   NOR2_X1 i_3417 (.A1(n_3841), .A2(n_3839), .ZN(n_3838));
   INV_X1 i_3418 (.A(n_3840), .ZN(n_3839));
   NAND3_X1 i_3419 (.A1(inputB[11]), .A2(inputA[14]), .A3(n_4032), .ZN(n_3840));
   AOI22_X1 i_3420 (.A1(inputB[10]), .A2(inputA[14]), .B1(inputB[11]), .B2(
      inputA[13]), .ZN(n_3841));
   INV_X1 i_3421 (.A(n_3842), .ZN(n_2433));
   AOI21_X1 i_3422 (.A(n_2430), .B1(n_2429), .B2(n_3952), .ZN(n_3842));
   INV_X1 i_3423 (.A(n_3843), .ZN(n_2423));
   AOI21_X1 i_3424 (.A(n_2420), .B1(n_2419), .B2(n_3957), .ZN(n_3843));
   XNOR2_X1 i_3425 (.A(n_2540), .B(n_3845), .ZN(n_2542));
   INV_X1 i_3426 (.A(n_3845), .ZN(n_3844));
   AOI21_X1 i_3427 (.A(n_2405), .B1(n_2404), .B2(n_3958), .ZN(n_3845));
   INV_X1 i_3428 (.A(n_3846), .ZN(n_2418));
   AOI21_X1 i_3429 (.A(n_2415), .B1(n_2414), .B2(n_3982), .ZN(n_3846));
   XOR2_X1 i_3430 (.A(n_2535), .B(n_3847), .Z(n_2537));
   XOR2_X1 i_3431 (.A(n_2515), .B(n_3850), .Z(n_3847));
   OAI21_X1 i_3432 (.A(n_3968), .B1(n_3973), .B2(n_3962), .ZN(n_3850));
   XOR2_X1 i_3433 (.A(n_2530), .B(n_3851), .Z(n_2532));
   XOR2_X1 i_3434 (.A(n_3853), .B(n_3852), .Z(n_3851));
   NAND2_X1 i_3435 (.A1(inputB[21]), .A2(inputA[3]), .ZN(n_3852));
   NAND2_X1 i_3436 (.A1(n_3857), .A2(n_3854), .ZN(n_3853));
   NAND3_X1 i_3437 (.A1(inputB[20]), .A2(inputA[5]), .A3(n_4018), .ZN(n_3854));
   INV_X1 i_3438 (.A(n_3858), .ZN(n_3857));
   AOI22_X1 i_3439 (.A1(inputB[19]), .A2(inputA[5]), .B1(inputB[20]), .B2(
      inputA[4]), .ZN(n_3858));
   INV_X1 i_3440 (.A(n_3859), .ZN(n_2413));
   AOI21_X1 i_3441 (.A(n_2410), .B1(n_2409), .B2(n_3976), .ZN(n_3859));
   INV_X1 i_3443 (.A(n_3860), .ZN(n_2398));
   AOI21_X1 i_3444 (.A(n_2395), .B1(n_2394), .B2(n_3988), .ZN(n_3860));
   INV_X1 i_3445 (.A(n_3861), .ZN(n_2403));
   AOI21_X1 i_3447 (.A(n_2400), .B1(n_2399), .B2(n_3996), .ZN(n_3861));
   XOR2_X1 i_3448 (.A(n_3863), .B(n_3862), .Z(n_2504));
   AND2_X1 i_3449 (.A1(inputB[0]), .A2(inputA[24]), .ZN(n_3862));
   AOI21_X1 i_3451 (.A(n_3864), .B1(n_3866), .B2(n_3865), .ZN(n_3863));
   NOR2_X1 i_3452 (.A1(n_3866), .A2(n_3865), .ZN(n_3864));
   AOI21_X1 i_3453 (.A(n_4045), .B1(n_4041), .B2(n_4039), .ZN(n_3865));
   INV_X1 i_3455 (.A(n_3867), .ZN(n_3866));
   OAI21_X1 i_3456 (.A(n_3993), .B1(n_3992), .B2(n_3989), .ZN(n_3867));
   XOR2_X1 i_3457 (.A(n_2510), .B(n_3868), .Z(n_2512));
   OAI21_X1 i_3459 (.A(n_4003), .B1(n_4000), .B2(n_3997), .ZN(n_3868));
   INV_X1 i_3460 (.A(n_3871), .ZN(n_2393));
   AOI21_X1 i_3461 (.A(n_2390), .B1(n_2389), .B2(n_3984), .ZN(n_3871));
   XOR2_X1 i_3463 (.A(n_3873), .B(n_3872), .Z(n_2448));
   NAND2_X1 i_3464 (.A1(inputB[24]), .A2(inputA[0]), .ZN(n_3872));
   NAND2_X1 i_3465 (.A1(n_3875), .A2(n_3874), .ZN(n_3873));
   NAND4_X1 i_3467 (.A1(inputB[22]), .A2(inputA[2]), .A3(inputB[23]), .A4(
      inputA[1]), .ZN(n_3874));
   INV_X1 i_3468 (.A(n_3878), .ZN(n_3875));
   AOI22_X1 i_3469 (.A1(inputB[22]), .A2(inputA[2]), .B1(inputB[23]), .B2(
      inputA[1]), .ZN(n_3878));
   XOR2_X1 i_3471 (.A(n_3880), .B(n_3879), .Z(n_2462));
   NAND2_X1 i_3472 (.A1(inputB[18]), .A2(inputA[6]), .ZN(n_3879));
   NAND2_X1 i_3473 (.A1(n_3882), .A2(n_3881), .ZN(n_3880));
   NAND4_X1 i_3475 (.A1(inputB[16]), .A2(inputA[8]), .A3(inputB[17]), .A4(
      inputA[7]), .ZN(n_3881));
   INV_X1 i_3476 (.A(n_3883), .ZN(n_3882));
   AOI22_X1 i_3477 (.A1(inputB[16]), .A2(inputA[8]), .B1(inputB[17]), .B2(
      inputA[7]), .ZN(n_3883));
   XOR2_X1 i_3479 (.A(n_3885), .B(n_3884), .Z(n_2469));
   NAND2_X1 i_3480 (.A1(inputB[15]), .A2(inputA[9]), .ZN(n_3884));
   NAND2_X1 i_3481 (.A1(n_3887), .A2(n_3886), .ZN(n_3885));
   NAND3_X1 i_3483 (.A1(inputB[14]), .A2(inputA[10]), .A3(n_4004), .ZN(n_3886));
   INV_X1 i_3484 (.A(n_3888), .ZN(n_3887));
   AOI21_X1 i_3485 (.A(n_4004), .B1(inputB[14]), .B2(inputA[10]), .ZN(n_3888));
   XOR2_X1 i_3487 (.A(n_3893), .B(n_3892), .Z(n_2483));
   NAND2_X1 i_3488 (.A1(inputB[9]), .A2(inputA[15]), .ZN(n_3892));
   NAND2_X1 i_3489 (.A1(n_3907), .A2(n_3896), .ZN(n_3893));
   NAND3_X1 i_3491 (.A1(inputB[7]), .A2(inputA[16]), .A3(n_3897), .ZN(n_3896));
   INV_X1 i_3492 (.A(n_3902), .ZN(n_3897));
   NAND2_X1 i_3493 (.A1(inputB[8]), .A2(inputA[17]), .ZN(n_3902));
   INV_X1 i_3495 (.A(n_3911), .ZN(n_3907));
   AOI22_X1 i_3496 (.A1(inputB[7]), .A2(inputA[17]), .B1(inputB[8]), .B2(
      inputA[16]), .ZN(n_3911));
   XOR2_X1 i_3497 (.A(n_3913), .B(n_3912), .Z(n_2490));
   NAND2_X1 i_3499 (.A1(inputB[6]), .A2(inputA[18]), .ZN(n_3912));
   OAI21_X1 i_3500 (.A(n_3916), .B1(n_3994), .B2(n_3917), .ZN(n_3913));
   NAND2_X1 i_3501 (.A1(n_3994), .A2(n_3917), .ZN(n_3916));
   INV_X1 i_3503 (.A(n_3922), .ZN(n_3917));
   NAND2_X1 i_3504 (.A1(inputB[5]), .A2(inputA[19]), .ZN(n_3922));
   INV_X1 i_3505 (.A(n_3927), .ZN(n_2383));
   AOI21_X1 i_3507 (.A(n_2380), .B1(n_2379), .B2(n_4011), .ZN(n_3927));
   INV_X1 i_3508 (.A(n_3928), .ZN(n_2388));
   AOI21_X1 i_3509 (.A(n_2385), .B1(n_2384), .B2(n_4012), .ZN(n_3928));
   OAI21_X1 i_3511 (.A(n_4015), .B1(n_4017), .B2(n_4013), .ZN(n_2333));
   OAI21_X1 i_3512 (.A(n_4021), .B1(n_4025), .B2(n_4019), .ZN(n_2340));
   NAND2_X1 i_3513 (.A1(n_4031), .A2(n_3932), .ZN(n_2354));
   NAND2_X1 i_3515 (.A1(n_4028), .A2(n_4026), .ZN(n_3932));
   OAI21_X1 i_3516 (.A(n_4036), .B1(n_4038), .B2(n_4034), .ZN(n_2361));
   XOR2_X1 i_3517 (.A(n_2439), .B(n_3933), .Z(n_2441));
   XOR2_X1 i_3518 (.A(n_2434), .B(n_3936), .Z(n_3933));
   XNOR2_X1 i_3519 (.A(n_2424), .B(n_3942), .ZN(n_3936));
   INV_X1 i_3520 (.A(n_3942), .ZN(n_3937));
   AOI21_X1 i_3521 (.A(n_2297), .B1(n_2296), .B2(n_4069), .ZN(n_3942));
   INV_X1 i_3522 (.A(n_3943), .ZN(n_2320));
   AOI21_X1 i_3523 (.A(n_2317), .B1(n_2316), .B2(n_4048), .ZN(n_3943));
   INV_X1 i_3524 (.A(n_3947), .ZN(n_2315));
   AOI21_X1 i_3525 (.A(n_2312), .B1(n_2311), .B2(n_4049), .ZN(n_3947));
   XNOR2_X1 i_3526 (.A(n_2429), .B(n_3953), .ZN(n_2431));
   INV_X1 i_3527 (.A(n_3953), .ZN(n_3952));
   AOI21_X1 i_3528 (.A(n_2302), .B1(n_2301), .B2(n_4052), .ZN(n_3953));
   INV_X1 i_3529 (.A(n_3956), .ZN(n_2310));
   AOI21_X1 i_3530 (.A(n_2307), .B1(n_2306), .B2(n_4064), .ZN(n_3956));
   XOR2_X1 i_3531 (.A(n_2419), .B(n_3957), .Z(n_2421));
   XOR2_X1 i_3532 (.A(n_2404), .B(n_3958), .Z(n_3957));
   XOR2_X1 i_3533 (.A(n_3967), .B(n_3962), .Z(n_3958));
   NAND2_X1 i_3534 (.A1(inputB[23]), .A2(inputA[0]), .ZN(n_3962));
   NAND2_X1 i_3535 (.A1(n_3972), .A2(n_3968), .ZN(n_3967));
   NAND4_X1 i_3536 (.A1(inputB[21]), .A2(inputA[2]), .A3(inputB[22]), .A4(
      inputA[1]), .ZN(n_3968));
   INV_X1 i_3537 (.A(n_3973), .ZN(n_3972));
   AOI22_X1 i_3538 (.A1(inputB[21]), .A2(inputA[2]), .B1(inputB[22]), .B2(
      inputA[1]), .ZN(n_3973));
   XNOR2_X1 i_3539 (.A(n_2409), .B(n_3977), .ZN(n_2411));
   INV_X1 i_3540 (.A(n_3977), .ZN(n_3976));
   AOI21_X1 i_3541 (.A(n_2282), .B1(n_2281), .B2(n_4110), .ZN(n_3977));
   XOR2_X1 i_3542 (.A(n_2414), .B(n_3982), .Z(n_2416));
   XNOR2_X1 i_3543 (.A(n_2389), .B(n_3987), .ZN(n_3982));
   INV_X1 i_3544 (.A(n_3987), .ZN(n_3984));
   AOI21_X1 i_3545 (.A(n_2262), .B1(n_2261), .B2(n_4152), .ZN(n_3987));
   XOR2_X1 i_3546 (.A(n_2394), .B(n_3988), .Z(n_2396));
   XOR2_X1 i_3547 (.A(n_3990), .B(n_3989), .Z(n_3988));
   NAND2_X1 i_3548 (.A1(inputB[5]), .A2(inputA[18]), .ZN(n_3989));
   NAND2_X1 i_3549 (.A1(n_3993), .A2(n_3991), .ZN(n_3990));
   INV_X1 i_3550 (.A(n_3992), .ZN(n_3991));
   AOI22_X1 i_3551 (.A1(inputB[3]), .A2(inputA[20]), .B1(inputB[4]), .B2(
      inputA[19]), .ZN(n_3992));
   NAND2_X1 i_3552 (.A1(n_4186), .A2(n_3994), .ZN(n_3993));
   INV_X1 i_3553 (.A(n_3995), .ZN(n_3994));
   NAND2_X1 i_3554 (.A1(inputB[4]), .A2(inputA[20]), .ZN(n_3995));
   XOR2_X1 i_3555 (.A(n_2399), .B(n_3996), .Z(n_2401));
   XOR2_X1 i_3556 (.A(n_3998), .B(n_3997), .Z(n_3996));
   NAND2_X1 i_3557 (.A1(inputB[14]), .A2(inputA[9]), .ZN(n_3997));
   NAND2_X1 i_3558 (.A1(n_4003), .A2(n_3999), .ZN(n_3998));
   INV_X1 i_3559 (.A(n_4000), .ZN(n_3999));
   AOI22_X1 i_3560 (.A1(inputB[12]), .A2(inputA[11]), .B1(inputB[13]), .B2(
      inputA[10]), .ZN(n_4000));
   NAND2_X1 i_3561 (.A1(n_4173), .A2(n_4004), .ZN(n_4003));
   AND2_X1 i_3562 (.A1(inputB[13]), .A2(inputA[11]), .ZN(n_4004));
   INV_X1 i_3563 (.A(n_4005), .ZN(n_2290));
   AOI21_X1 i_3564 (.A(n_2287), .B1(n_2286), .B2(n_4053), .ZN(n_4005));
   INV_X1 i_3565 (.A(n_4006), .ZN(n_2295));
   AOI21_X1 i_3566 (.A(n_2292), .B1(n_2291), .B2(n_4075), .ZN(n_4006));
   INV_X1 i_3567 (.A(n_4007), .ZN(n_2275));
   AOI21_X1 i_3568 (.A(n_2272), .B1(n_2271), .B2(n_4134), .ZN(n_4007));
   INV_X1 i_3569 (.A(n_4010), .ZN(n_2280));
   AOI21_X1 i_3570 (.A(n_2277), .B1(n_2276), .B2(n_4080), .ZN(n_4010));
   XOR2_X1 i_3571 (.A(n_2379), .B(n_4011), .Z(n_2381));
   AOI21_X1 i_3572 (.A(n_4099), .B1(n_4104), .B2(n_4084), .ZN(n_4011));
   XOR2_X1 i_3573 (.A(n_2384), .B(n_4012), .Z(n_2386));
   OAI21_X1 i_3574 (.A(n_4119), .B1(n_4129), .B2(n_4114), .ZN(n_4012));
   XOR2_X1 i_3575 (.A(n_4014), .B(n_4013), .Z(n_2332));
   NAND2_X1 i_3576 (.A1(inputB[20]), .A2(inputA[3]), .ZN(n_4013));
   NAND2_X1 i_3577 (.A1(n_4016), .A2(n_4015), .ZN(n_4014));
   NAND3_X1 i_3578 (.A1(inputB[18]), .A2(inputA[5]), .A3(n_4018), .ZN(n_4015));
   INV_X1 i_3579 (.A(n_4017), .ZN(n_4016));
   AOI21_X1 i_3580 (.A(n_4018), .B1(inputB[18]), .B2(inputA[5]), .ZN(n_4017));
   AND2_X1 i_3581 (.A1(inputB[19]), .A2(inputA[4]), .ZN(n_4018));
   XOR2_X1 i_3582 (.A(n_4020), .B(n_4019), .Z(n_2339));
   NAND2_X1 i_3583 (.A1(inputB[17]), .A2(inputA[6]), .ZN(n_4019));
   NAND2_X1 i_3584 (.A1(n_4024), .A2(n_4021), .ZN(n_4020));
   NAND4_X1 i_3585 (.A1(inputB[15]), .A2(inputA[8]), .A3(inputB[16]), .A4(
      inputA[7]), .ZN(n_4021));
   INV_X1 i_3586 (.A(n_4025), .ZN(n_4024));
   AOI22_X1 i_3587 (.A1(inputB[15]), .A2(inputA[8]), .B1(inputB[16]), .B2(
      inputA[7]), .ZN(n_4025));
   XOR2_X1 i_3588 (.A(n_4027), .B(n_4026), .Z(n_2353));
   AND2_X1 i_3589 (.A1(inputB[11]), .A2(inputA[12]), .ZN(n_4026));
   AND2_X1 i_3591 (.A1(n_4031), .A2(n_4028), .ZN(n_4027));
   NAND2_X1 i_3592 (.A1(n_4109), .A2(n_4033), .ZN(n_4028));
   NAND2_X1 i_3593 (.A1(n_4105), .A2(n_4032), .ZN(n_4031));
   INV_X1 i_3595 (.A(n_4033), .ZN(n_4032));
   NAND2_X1 i_3596 (.A1(inputB[10]), .A2(inputA[13]), .ZN(n_4033));
   XOR2_X1 i_3597 (.A(n_4035), .B(n_4034), .Z(n_2360));
   NAND2_X1 i_3599 (.A1(inputB[8]), .A2(inputA[15]), .ZN(n_4034));
   NAND2_X1 i_3600 (.A1(n_4037), .A2(n_4036), .ZN(n_4035));
   NAND3_X1 i_3601 (.A1(inputB[7]), .A2(inputA[17]), .A3(n_4179), .ZN(n_4036));
   INV_X1 i_3603 (.A(n_4038), .ZN(n_4037));
   AOI22_X1 i_3604 (.A1(inputB[6]), .A2(inputA[17]), .B1(inputB[7]), .B2(
      inputA[16]), .ZN(n_4038));
   XOR2_X1 i_3605 (.A(n_4040), .B(n_4039), .Z(n_2374));
   AND2_X1 i_3607 (.A1(inputB[2]), .A2(inputA[21]), .ZN(n_4039));
   NOR2_X1 i_3608 (.A1(n_4045), .A2(n_4042), .ZN(n_4040));
   INV_X1 i_3609 (.A(n_4042), .ZN(n_4041));
   AOI21_X1 i_3611 (.A(n_4146), .B1(inputB[0]), .B2(inputA[23]), .ZN(n_4042));
   AND3_X1 i_3612 (.A1(inputB[0]), .A2(inputA[23]), .A3(n_4146), .ZN(n_4045));
   INV_X1 i_3613 (.A(n_4046), .ZN(n_2270));
   AOI21_X1 i_3615 (.A(n_2267), .B1(n_2266), .B2(n_4054), .ZN(n_4046));
   OAI21_X1 i_3616 (.A(n_4158), .B1(n_4160), .B2(n_4154), .ZN(n_2207));
   OAI21_X1 i_3617 (.A(n_4163), .B1(n_4166), .B2(n_4161), .ZN(n_2221));
   OAI21_X1 i_3619 (.A(n_4169), .B1(n_4172), .B2(n_4167), .ZN(n_2228));
   AOI22_X1 i_3620 (.A1(n_4203), .A2(n_4180), .B1(n_4176), .B2(n_4174), .ZN(
      n_2242));
   NAND2_X1 i_3621 (.A1(n_4184), .A2(n_4047), .ZN(n_2249));
   NAND2_X1 i_3623 (.A1(n_4183), .A2(n_4181), .ZN(n_4047));
   XOR2_X1 i_3624 (.A(n_2316), .B(n_4048), .Z(n_2318));
   XOR2_X1 i_3625 (.A(n_2311), .B(n_4049), .Z(n_4048));
   XOR2_X1 i_3627 (.A(n_2301), .B(n_4052), .Z(n_4049));
   XOR2_X1 i_3628 (.A(n_2286), .B(n_4053), .Z(n_4052));
   XOR2_X1 i_3629 (.A(n_2266), .B(n_4054), .Z(n_4053));
   OAI21_X1 i_3631 (.A(n_4304), .B1(n_4306), .B2(n_4301), .ZN(n_4054));
   INV_X1 i_3632 (.A(n_4055), .ZN(n_2201));
   AOI21_X1 i_3633 (.A(n_2198), .B1(n_2197), .B2(n_4190), .ZN(n_4055));
   INV_X1 i_3635 (.A(n_4059), .ZN(n_2196));
   AOI21_X1 i_3636 (.A(n_2193), .B1(n_2192), .B2(n_4192), .ZN(n_4059));
   XNOR2_X1 i_3637 (.A(n_2306), .B(n_4065), .ZN(n_2308));
   INV_X1 i_3639 (.A(n_4065), .ZN(n_4064));
   AOI21_X1 i_3640 (.A(n_2183), .B1(n_2182), .B2(n_4193), .ZN(n_4065));
   INV_X1 i_3641 (.A(n_4068), .ZN(n_2191));
   AOI21_X1 i_3643 (.A(n_2188), .B1(n_2187), .B2(n_4207), .ZN(n_4068));
   XNOR2_X1 i_3644 (.A(n_2296), .B(n_4074), .ZN(n_2298));
   INV_X1 i_3645 (.A(n_4074), .ZN(n_4069));
   AOI21_X1 i_3647 (.A(n_2168), .B1(n_2167), .B2(n_4268), .ZN(n_4074));
   XNOR2_X1 i_3648 (.A(n_2291), .B(n_4078), .ZN(n_2293));
   INV_X1 i_3649 (.A(n_4078), .ZN(n_4075));
   AOI21_X1 i_3651 (.A(n_2158), .B1(n_2157), .B2(n_4194), .ZN(n_4078));
   INV_X1 i_3652 (.A(n_4079), .ZN(n_2181));
   AOI21_X1 i_3653 (.A(n_2178), .B1(n_2177), .B2(n_4238), .ZN(n_4079));
   XOR2_X1 i_3655 (.A(n_2276), .B(n_4080), .Z(n_2278));
   XOR2_X1 i_3656 (.A(n_4089), .B(n_4084), .Z(n_4080));
   NAND2_X1 i_3657 (.A1(inputB[10]), .A2(inputA[12]), .ZN(n_4084));
   NAND2_X1 i_3659 (.A1(n_4104), .A2(n_4094), .ZN(n_4089));
   INV_X1 i_3660 (.A(n_4099), .ZN(n_4094));
   AOI22_X1 i_3661 (.A1(inputB[8]), .A2(inputA[14]), .B1(inputB[9]), .B2(
      inputA[13]), .ZN(n_4099));
   NAND2_X1 i_3663 (.A1(n_4324), .A2(n_4105), .ZN(n_4104));
   INV_X1 i_3664 (.A(n_4109), .ZN(n_4105));
   NAND2_X1 i_3665 (.A1(inputB[9]), .A2(inputA[14]), .ZN(n_4109));
   XOR2_X1 i_3666 (.A(n_2281), .B(n_4110), .Z(n_2283));
   XOR2_X1 i_3667 (.A(n_4115), .B(n_4114), .Z(n_4110));
   NAND2_X1 i_3668 (.A1(inputB[19]), .A2(inputA[3]), .ZN(n_4114));
   NAND2_X1 i_3669 (.A1(n_4124), .A2(n_4119), .ZN(n_4115));
   NAND3_X1 i_3670 (.A1(inputB[18]), .A2(inputA[4]), .A3(n_4312), .ZN(n_4119));
   INV_X1 i_3671 (.A(n_4129), .ZN(n_4124));
   AOI21_X1 i_3672 (.A(n_4312), .B1(inputB[18]), .B2(inputA[4]), .ZN(n_4129));
   INV_X1 i_3673 (.A(n_4130), .ZN(n_2176));
   AOI21_X1 i_3674 (.A(n_2173), .B1(n_2172), .B2(n_4208), .ZN(n_4130));
   XOR2_X1 i_3675 (.A(n_2271), .B(n_4134), .Z(n_2273));
   AOI21_X1 i_3676 (.A(n_4138), .B1(n_4149), .B2(n_4148), .ZN(n_4134));
   INV_X1 i_3677 (.A(n_4139), .ZN(n_4138));
   OAI21_X1 i_3678 (.A(n_2255), .B1(n_4149), .B2(n_4144), .ZN(n_4139));
   AOI21_X1 i_3679 (.A(n_4148), .B1(n_4149), .B2(n_4144), .ZN(n_2255));
   NAND2_X1 i_3680 (.A1(n_4283), .A2(n_4146), .ZN(n_4144));
   AND2_X1 i_3681 (.A1(inputB[1]), .A2(inputA[22]), .ZN(n_4146));
   AOI22_X1 i_3682 (.A1(inputB[0]), .A2(inputA[22]), .B1(inputB[1]), .B2(
      inputA[21]), .ZN(n_4148));
   INV_X1 i_3683 (.A(n_4150), .ZN(n_4149));
   AOI21_X1 i_3684 (.A(n_4330), .B1(n_4333), .B2(n_4327), .ZN(n_4150));
   INV_X1 i_3685 (.A(n_4151), .ZN(n_2166));
   AOI21_X1 i_3686 (.A(n_2163), .B1(n_2162), .B2(n_4247), .ZN(n_4151));
   XOR2_X1 i_3687 (.A(n_2261), .B(n_4152), .Z(n_2263));
   OAI21_X1 i_3688 (.A(n_4318), .B1(n_4320), .B2(n_4315), .ZN(n_4152));
   INV_X1 i_3689 (.A(n_4153), .ZN(n_2156));
   AOI21_X1 i_3690 (.A(n_2153), .B1(n_2152), .B2(n_4269), .ZN(n_4153));
   XOR2_X1 i_3691 (.A(n_4155), .B(n_4154), .Z(n_2206));
   NAND2_X1 i_3692 (.A1(inputB[22]), .A2(inputA[0]), .ZN(n_4154));
   NAND2_X1 i_3693 (.A1(n_4159), .A2(n_4158), .ZN(n_4155));
   NAND4_X1 i_3694 (.A1(inputB[20]), .A2(inputA[2]), .A3(inputB[21]), .A4(
      inputA[1]), .ZN(n_4158));
   INV_X1 i_3695 (.A(n_4160), .ZN(n_4159));
   AOI22_X1 i_3696 (.A1(inputB[20]), .A2(inputA[2]), .B1(inputB[21]), .B2(
      inputA[1]), .ZN(n_4160));
   XOR2_X1 i_3697 (.A(n_4162), .B(n_4161), .Z(n_2220));
   NAND2_X1 i_3698 (.A1(inputB[16]), .A2(inputA[6]), .ZN(n_4161));
   NAND2_X1 i_3699 (.A1(n_4165), .A2(n_4163), .ZN(n_4162));
   NAND3_X1 i_3700 (.A1(inputB[15]), .A2(inputA[7]), .A3(n_4264), .ZN(n_4163));
   INV_X1 i_3701 (.A(n_4166), .ZN(n_4165));
   AOI21_X1 i_3702 (.A(n_4264), .B1(inputB[15]), .B2(inputA[7]), .ZN(n_4166));
   XOR2_X1 i_3703 (.A(n_4168), .B(n_4167), .Z(n_2227));
   NAND2_X1 i_3704 (.A1(inputB[13]), .A2(inputA[9]), .ZN(n_4167));
   NAND2_X1 i_3705 (.A1(n_4171), .A2(n_4169), .ZN(n_4168));
   NAND3_X1 i_3706 (.A1(inputB[11]), .A2(inputA[11]), .A3(n_4173), .ZN(n_4169));
   INV_X1 i_3707 (.A(n_4172), .ZN(n_4171));
   AOI21_X1 i_3708 (.A(n_4173), .B1(inputB[11]), .B2(inputA[11]), .ZN(n_4172));
   AND2_X1 i_3709 (.A1(inputB[12]), .A2(inputA[10]), .ZN(n_4173));
   XOR2_X1 i_3710 (.A(n_4175), .B(n_4174), .Z(n_2241));
   NAND2_X1 i_3711 (.A1(inputB[7]), .A2(inputA[15]), .ZN(n_4174));
   OAI21_X1 i_3712 (.A(n_4176), .B1(n_4202), .B2(n_4179), .ZN(n_4175));
   NAND2_X1 i_3713 (.A1(n_4202), .A2(n_4179), .ZN(n_4176));
   INV_X1 i_3714 (.A(n_4180), .ZN(n_4179));
   NAND2_X1 i_3715 (.A1(inputB[6]), .A2(inputA[16]), .ZN(n_4180));
   XOR2_X1 i_3716 (.A(n_4182), .B(n_4181), .Z(n_2248));
   AND2_X1 i_3717 (.A1(inputB[4]), .A2(inputA[18]), .ZN(n_4181));
   AND2_X1 i_3718 (.A1(n_4184), .A2(n_4183), .ZN(n_4182));
   NAND2_X1 i_3719 (.A1(n_4335), .A2(n_4187), .ZN(n_4183));
   NAND2_X1 i_3720 (.A1(n_4334), .A2(n_4186), .ZN(n_4184));
   INV_X1 i_3721 (.A(n_4187), .ZN(n_4186));
   NAND2_X1 i_3722 (.A1(inputB[3]), .A2(inputA[19]), .ZN(n_4187));
   AOI21_X1 i_3723 (.A(n_4188), .B1(n_4292), .B2(n_4289), .ZN(n_2142));
   NOR2_X1 i_3724 (.A1(n_4288), .A2(n_4283), .ZN(n_4188));
   INV_X1 i_3725 (.A(n_4189), .ZN(n_2151));
   AOI21_X1 i_3726 (.A(n_2148), .B1(n_2147), .B2(n_4298), .ZN(n_4189));
   OAI21_X1 i_3727 (.A(n_4309), .B1(n_4314), .B2(n_4307), .ZN(n_2100));
   OAI21_X1 i_3728 (.A(n_4263), .B1(n_4262), .B2(n_4248), .ZN(n_2107));
   AOI22_X1 i_3729 (.A1(n_4438), .A2(n_4326), .B1(n_4323), .B2(n_4321), .ZN(
      n_2121));
   OAI21_X1 i_3730 (.A(n_4201), .B1(n_4200), .B2(n_4195), .ZN(n_2128));
   XOR2_X1 i_3731 (.A(n_2197), .B(n_4190), .Z(n_2199));
   XOR2_X1 i_3732 (.A(n_2192), .B(n_4192), .Z(n_4190));
   XOR2_X1 i_3733 (.A(n_2182), .B(n_4193), .Z(n_4192));
   XOR2_X1 i_3734 (.A(n_2157), .B(n_4194), .Z(n_4193));
   XOR2_X1 i_3735 (.A(n_4196), .B(n_4195), .Z(n_4194));
   NAND2_X1 i_3736 (.A1(inputB[6]), .A2(inputA[15]), .ZN(n_4195));
   NAND2_X1 i_3737 (.A1(n_4201), .A2(n_4197), .ZN(n_4196));
   INV_X1 i_3739 (.A(n_4200), .ZN(n_4197));
   AOI22_X1 i_3740 (.A1(inputB[4]), .A2(inputA[17]), .B1(inputB[5]), .B2(
      inputA[16]), .ZN(n_4200));
   NAND2_X1 i_3741 (.A1(n_4452), .A2(n_4202), .ZN(n_4201));
   INV_X1 i_3743 (.A(n_4203), .ZN(n_4202));
   NAND2_X1 i_3744 (.A1(inputB[5]), .A2(inputA[17]), .ZN(n_4203));
   INV_X1 i_3745 (.A(n_4204), .ZN(n_2087));
   AOI21_X1 i_3747 (.A(n_2084), .B1(n_2083), .B2(n_4205), .ZN(n_4204));
   XOR2_X1 i_3748 (.A(n_2078), .B(n_4213), .Z(n_4205));
   XOR2_X1 i_3749 (.A(n_2187), .B(n_4207), .Z(n_2189));
   XNOR2_X1 i_3751 (.A(n_2172), .B(n_4209), .ZN(n_4207));
   INV_X1 i_3752 (.A(n_4209), .ZN(n_4208));
   AOI21_X1 i_3753 (.A(n_2054), .B1(n_2053), .B2(n_4228), .ZN(n_4209));
   INV_X1 i_3755 (.A(n_4212), .ZN(n_2082));
   AOI21_X1 i_3756 (.A(n_2079), .B1(n_2078), .B2(n_4213), .ZN(n_4212));
   XOR2_X1 i_3757 (.A(n_2068), .B(n_4223), .Z(n_4213));
   INV_X1 i_3759 (.A(n_4214), .ZN(n_2077));
   AOI21_X1 i_3760 (.A(n_2074), .B1(n_2073), .B2(n_4343), .ZN(n_4214));
   INV_X1 i_3761 (.A(n_4218), .ZN(n_2072));
   AOI21_X1 i_3763 (.A(n_2069), .B1(n_2068), .B2(n_4223), .ZN(n_4218));
   XOR2_X1 i_3764 (.A(n_2053), .B(n_4228), .Z(n_4223));
   XNOR2_X1 i_3765 (.A(n_4337), .B(n_4233), .ZN(n_4228));
   AOI21_X1 i_3767 (.A(n_4341), .B1(n_4504), .B2(n_4340), .ZN(n_4233));
   XNOR2_X1 i_3768 (.A(n_2177), .B(n_4239), .ZN(n_2179));
   INV_X1 i_3769 (.A(n_4239), .ZN(n_4238));
   AOI21_X1 i_3771 (.A(n_2059), .B1(n_2058), .B2(n_4344), .ZN(n_4239));
   INV_X1 i_3772 (.A(n_4243), .ZN(n_2067));
   AOI21_X1 i_3773 (.A(n_2064), .B1(n_2063), .B2(n_4350), .ZN(n_4243));
   XOR2_X1 i_3775 (.A(n_2162), .B(n_4247), .Z(n_2164));
   XOR2_X1 i_3776 (.A(n_4253), .B(n_4248), .Z(n_4247));
   NAND2_X1 i_3777 (.A1(inputB[15]), .A2(inputA[6]), .ZN(n_4248));
   NAND2_X1 i_3779 (.A1(n_4263), .A2(n_4258), .ZN(n_4253));
   INV_X1 i_3780 (.A(n_4262), .ZN(n_4258));
   AOI22_X1 i_3781 (.A1(inputB[13]), .A2(inputA[8]), .B1(inputB[14]), .B2(
      inputA[7]), .ZN(n_4262));
   NAND2_X1 i_3783 (.A1(n_4417), .A2(n_4264), .ZN(n_4263));
   AND2_X1 i_3784 (.A1(inputB[14]), .A2(inputA[8]), .ZN(n_4264));
   XOR2_X1 i_3785 (.A(n_2167), .B(n_4268), .Z(n_2169));
   XNOR2_X1 i_3787 (.A(n_2152), .B(n_4273), .ZN(n_4268));
   INV_X1 i_3788 (.A(n_4273), .ZN(n_4269));
   AOI21_X1 i_3789 (.A(n_2039), .B1(n_2038), .B2(n_4383), .ZN(n_4273));
   INV_X1 i_3791 (.A(n_4278), .ZN(n_2047));
   AOI21_X1 i_3792 (.A(n_2044), .B1(n_2043), .B2(n_4351), .ZN(n_4278));
   INV_X1 i_3793 (.A(n_4282), .ZN(n_2052));
   AOI21_X1 i_3795 (.A(n_2049), .B1(n_2048), .B2(n_4360), .ZN(n_4282));
   XOR2_X1 i_3796 (.A(n_4284), .B(n_4283), .Z(n_2141));
   AND2_X1 i_3797 (.A1(inputB[0]), .A2(inputA[21]), .ZN(n_4283));
   AOI21_X1 i_3799 (.A(n_4288), .B1(n_4292), .B2(n_4289), .ZN(n_4284));
   NOR2_X1 i_3800 (.A1(n_4292), .A2(n_4289), .ZN(n_4288));
   AOI22_X1 i_3801 (.A1(n_4479), .A2(n_4452), .B1(n_4450), .B2(n_4443), .ZN(
      n_4289));
   INV_X1 i_3803 (.A(n_4293), .ZN(n_4292));
   OAI21_X1 i_3804 (.A(n_4356), .B1(n_4359), .B2(n_4354), .ZN(n_4293));
   XOR2_X1 i_3805 (.A(n_2147), .B(n_4298), .Z(n_2149));
   NAND2_X1 i_3807 (.A1(n_4413), .A2(n_4300), .ZN(n_4298));
   NAND2_X1 i_3808 (.A1(n_4408), .A2(n_4403), .ZN(n_4300));
   XOR2_X1 i_3809 (.A(n_4303), .B(n_4301), .Z(n_2092));
   NAND2_X1 i_3810 (.A1(inputB[21]), .A2(inputA[0]), .ZN(n_4301));
   NAND2_X1 i_3811 (.A1(n_4305), .A2(n_4304), .ZN(n_4303));
   NAND3_X1 i_3812 (.A1(inputB[20]), .A2(inputA[1]), .A3(n_4340), .ZN(n_4304));
   INV_X1 i_3813 (.A(n_4306), .ZN(n_4305));
   AOI21_X1 i_3814 (.A(n_4340), .B1(inputB[20]), .B2(inputA[1]), .ZN(n_4306));
   XOR2_X1 i_3815 (.A(n_4308), .B(n_4307), .Z(n_2099));
   NAND2_X1 i_3816 (.A1(inputB[18]), .A2(inputA[3]), .ZN(n_4307));
   NAND2_X1 i_3817 (.A1(n_4313), .A2(n_4309), .ZN(n_4308));
   NAND3_X1 i_3818 (.A1(inputB[16]), .A2(inputA[4]), .A3(n_4312), .ZN(n_4309));
   AND2_X1 i_3819 (.A1(inputB[17]), .A2(inputA[5]), .ZN(n_4312));
   INV_X1 i_3820 (.A(n_4314), .ZN(n_4313));
   AOI22_X1 i_3821 (.A1(inputB[16]), .A2(inputA[5]), .B1(inputB[17]), .B2(
      inputA[4]), .ZN(n_4314));
   XOR2_X1 i_3822 (.A(n_4316), .B(n_4315), .Z(n_2113));
   NAND2_X1 i_3823 (.A1(inputB[12]), .A2(inputA[9]), .ZN(n_4315));
   NAND2_X1 i_3824 (.A1(n_4319), .A2(n_4318), .ZN(n_4316));
   NAND3_X1 i_3825 (.A1(inputB[11]), .A2(inputA[10]), .A3(n_4372), .ZN(n_4318));
   INV_X1 i_3826 (.A(n_4320), .ZN(n_4319));
   AOI21_X1 i_3827 (.A(n_4372), .B1(inputB[11]), .B2(inputA[10]), .ZN(n_4320));
   XOR2_X1 i_3828 (.A(n_4322), .B(n_4321), .Z(n_2120));
   NAND2_X1 i_3829 (.A1(inputB[9]), .A2(inputA[12]), .ZN(n_4321));
   OAI21_X1 i_3830 (.A(n_4323), .B1(n_4434), .B2(n_4324), .ZN(n_4322));
   NAND2_X1 i_3831 (.A1(n_4434), .A2(n_4324), .ZN(n_4323));
   INV_X1 i_3832 (.A(n_4326), .ZN(n_4324));
   NAND2_X1 i_3833 (.A1(inputB[8]), .A2(inputA[13]), .ZN(n_4326));
   XOR2_X1 i_3834 (.A(n_4328), .B(n_4327), .Z(n_2134));
   NAND2_X1 i_3835 (.A1(inputB[3]), .A2(inputA[18]), .ZN(n_4327));
   NAND2_X1 i_3836 (.A1(n_4333), .A2(n_4329), .ZN(n_4328));
   INV_X1 i_3837 (.A(n_4330), .ZN(n_4329));
   AOI22_X1 i_3838 (.A1(inputB[1]), .A2(inputA[20]), .B1(inputB[2]), .B2(
      inputA[19]), .ZN(n_4330));
   NAND2_X1 i_3839 (.A1(n_4543), .A2(n_4334), .ZN(n_4333));
   INV_X1 i_3840 (.A(n_4335), .ZN(n_4334));
   NAND2_X1 i_3841 (.A1(inputB[2]), .A2(inputA[20]), .ZN(n_4335));
   INV_X1 i_3842 (.A(n_4336), .ZN(n_2037));
   AOI21_X1 i_3843 (.A(n_2034), .B1(n_2033), .B2(n_4345), .ZN(n_4336));
   OAI21_X1 i_3844 (.A(n_4339), .B1(n_4341), .B2(n_4337), .ZN(n_1987));
   NAND2_X1 i_3845 (.A1(inputB[20]), .A2(inputA[0]), .ZN(n_4337));
   NAND2_X1 i_3846 (.A1(n_4504), .A2(n_4340), .ZN(n_4339));
   AND2_X1 i_3847 (.A1(inputB[19]), .A2(inputA[2]), .ZN(n_4340));
   AOI22_X1 i_3848 (.A1(inputB[18]), .A2(inputA[2]), .B1(inputB[19]), .B2(
      inputA[1]), .ZN(n_4341));
   OAI21_X1 i_3849 (.A(n_4393), .B1(n_4398), .B2(n_4388), .ZN(n_1994));
   OAI21_X1 i_3850 (.A(n_4368), .B1(n_4364), .B2(n_4361), .ZN(n_2008));
   OAI21_X1 i_3851 (.A(n_4433), .B1(n_4442), .B2(n_4423), .ZN(n_2015));
   INV_X1 i_3852 (.A(n_4342), .ZN(n_1981));
   AOI21_X1 i_3853 (.A(n_1978), .B1(n_1977), .B2(n_4456), .ZN(n_4342));
   XOR2_X1 i_3854 (.A(n_2073), .B(n_4343), .Z(n_2075));
   XOR2_X1 i_3855 (.A(n_2058), .B(n_4344), .Z(n_4343));
   XOR2_X1 i_3856 (.A(n_2033), .B(n_4345), .Z(n_4344));
   OAI21_X1 i_3857 (.A(n_4512), .B1(n_4514), .B2(n_4510), .ZN(n_4345));
   INV_X1 i_3858 (.A(n_4347), .ZN(n_1976));
   AOI21_X1 i_3859 (.A(n_1973), .B1(n_1972), .B2(n_4457), .ZN(n_4347));
   INV_X1 i_3860 (.A(n_4348), .ZN(n_1971));
   AOI21_X1 i_3861 (.A(n_1968), .B1(n_1967), .B2(n_4466), .ZN(n_4348));
   INV_X1 i_3862 (.A(n_4349), .ZN(n_1966));
   AOI21_X1 i_3863 (.A(n_1963), .B1(n_1962), .B2(n_4458), .ZN(n_4349));
   XOR2_X1 i_3864 (.A(n_2063), .B(n_4350), .Z(n_2065));
   XOR2_X1 i_3865 (.A(n_2043), .B(n_4351), .Z(n_4350));
   XOR2_X1 i_3866 (.A(n_4355), .B(n_4354), .Z(n_4351));
   NAND2_X1 i_3867 (.A1(inputB[2]), .A2(inputA[18]), .ZN(n_4354));
   NAND2_X1 i_3868 (.A1(n_4357), .A2(n_4356), .ZN(n_4355));
   NAND3_X1 i_3869 (.A1(inputB[0]), .A2(inputA[20]), .A3(n_4543), .ZN(n_4356));
   INV_X1 i_3870 (.A(n_4359), .ZN(n_4357));
   AOI21_X1 i_3871 (.A(n_4543), .B1(inputB[0]), .B2(inputA[20]), .ZN(n_4359));
   XOR2_X1 i_3872 (.A(n_2048), .B(n_4360), .Z(n_2050));
   XOR2_X1 i_3873 (.A(n_4362), .B(n_4361), .Z(n_4360));
   NAND2_X1 i_3875 (.A1(inputB[11]), .A2(inputA[9]), .ZN(n_4361));
   NAND2_X1 i_3876 (.A1(n_4368), .A2(n_4363), .ZN(n_4362));
   INV_X1 i_3877 (.A(n_4364), .ZN(n_4363));
   AOI22_X1 i_3879 (.A1(inputB[9]), .A2(inputA[11]), .B1(inputB[10]), .B2(
      inputA[10]), .ZN(n_4364));
   NAND2_X1 i_3880 (.A1(n_4517), .A2(n_4372), .ZN(n_4368));
   AND2_X1 i_3881 (.A1(inputB[10]), .A2(inputA[11]), .ZN(n_4372));
   INV_X1 i_3883 (.A(n_4373), .ZN(n_1956));
   AOI21_X1 i_3884 (.A(n_1953), .B1(n_1952), .B2(n_4459), .ZN(n_4373));
   INV_X1 i_3885 (.A(n_4378), .ZN(n_1961));
   AOI21_X1 i_3887 (.A(n_1958), .B1(n_1957), .B2(n_4470), .ZN(n_4378));
   INV_X1 i_3888 (.A(n_4379), .ZN(n_1946));
   AOI21_X1 i_3889 (.A(n_1943), .B1(n_1942), .B2(n_4472), .ZN(n_4379));
   INV_X1 i_3891 (.A(n_4382), .ZN(n_1951));
   AOI21_X1 i_3892 (.A(n_1948), .B1(n_1947), .B2(n_4483), .ZN(n_4382));
   XOR2_X1 i_3893 (.A(n_2038), .B(n_4383), .Z(n_2040));
   OAI21_X1 i_3895 (.A(n_4499), .B1(n_4501), .B2(n_4497), .ZN(n_4383));
   INV_X1 i_3896 (.A(n_4384), .ZN(n_1941));
   AOI21_X1 i_3897 (.A(n_1938), .B1(n_1937), .B2(n_4462), .ZN(n_4384));
   XOR2_X1 i_3899 (.A(n_4389), .B(n_4388), .Z(n_1993));
   NAND2_X1 i_3900 (.A1(inputB[17]), .A2(inputA[3]), .ZN(n_4388));
   NAND2_X1 i_3901 (.A1(n_4397), .A2(n_4393), .ZN(n_4389));
   NAND4_X1 i_3903 (.A1(inputB[15]), .A2(inputA[4]), .A3(inputB[16]), .A4(
      inputA[5]), .ZN(n_4393));
   INV_X1 i_3904 (.A(n_4398), .ZN(n_4397));
   AOI22_X1 i_3905 (.A1(inputB[15]), .A2(inputA[5]), .B1(inputB[16]), .B2(
      inputA[4]), .ZN(n_4398));
   XOR2_X1 i_3907 (.A(n_4404), .B(n_4403), .Z(n_2000));
   AND2_X1 i_3908 (.A1(inputB[14]), .A2(inputA[6]), .ZN(n_4403));
   AND2_X1 i_3909 (.A1(n_4413), .A2(n_4408), .ZN(n_4404));
   NAND2_X1 i_3911 (.A1(n_4488), .A2(n_4418), .ZN(n_4408));
   NAND2_X1 i_3912 (.A1(n_4487), .A2(n_4417), .ZN(n_4413));
   INV_X1 i_3913 (.A(n_4418), .ZN(n_4417));
   NAND2_X1 i_3915 (.A1(inputB[13]), .A2(inputA[7]), .ZN(n_4418));
   XOR2_X1 i_3916 (.A(n_4428), .B(n_4423), .Z(n_2014));
   NAND2_X1 i_3917 (.A1(inputB[8]), .A2(inputA[12]), .ZN(n_4423));
   NAND2_X1 i_3919 (.A1(n_4439), .A2(n_4433), .ZN(n_4428));
   NAND3_X1 i_3920 (.A1(inputB[6]), .A2(inputA[13]), .A3(n_4434), .ZN(n_4433));
   INV_X1 i_3921 (.A(n_4438), .ZN(n_4434));
   NAND2_X1 i_3923 (.A1(inputB[7]), .A2(inputA[14]), .ZN(n_4438));
   INV_X1 i_3924 (.A(n_4442), .ZN(n_4439));
   AOI22_X1 i_3925 (.A1(inputB[6]), .A2(inputA[14]), .B1(inputB[7]), .B2(
      inputA[13]), .ZN(n_4442));
   XOR2_X1 i_3927 (.A(n_4448), .B(n_4443), .Z(n_2021));
   AND2_X1 i_3928 (.A1(inputB[5]), .A2(inputA[15]), .ZN(n_4443));
   AOI22_X1 i_3929 (.A1(n_4479), .A2(n_4452), .B1(n_4480), .B2(n_4453), .ZN(
      n_4448));
   NAND2_X1 i_3931 (.A1(n_4480), .A2(n_4453), .ZN(n_4450));
   INV_X1 i_3932 (.A(n_4453), .ZN(n_4452));
   NAND2_X1 i_3933 (.A1(inputB[4]), .A2(inputA[16]), .ZN(n_4453));
   INV_X1 i_3935 (.A(n_4454), .ZN(n_1926));
   AOI22_X1 i_3936 (.A1(n_4614), .A2(n_4543), .B1(n_4537), .B2(n_4534), .ZN(
      n_4454));
   INV_X1 i_3937 (.A(n_4455), .ZN(n_1936));
   AOI21_X1 i_3939 (.A(n_1933), .B1(n_1932), .B2(n_4496), .ZN(n_4455));
   OAI21_X1 i_3940 (.A(n_4507), .B1(n_4509), .B2(n_4505), .ZN(n_1892));
   OAI21_X1 i_3941 (.A(n_4486), .B1(n_4491), .B2(n_4490), .ZN(n_1899));
   OAI21_X1 i_3943 (.A(n_4528), .B1(n_4533), .B2(n_4518), .ZN(n_1913));
   OAI21_X1 i_3944 (.A(n_4478), .B1(n_4477), .B2(n_4473), .ZN(n_1920));
   XOR2_X1 i_3945 (.A(n_1977), .B(n_4456), .Z(n_1979));
   XOR2_X1 i_3946 (.A(n_1972), .B(n_4457), .Z(n_4456));
   XOR2_X1 i_3947 (.A(n_1962), .B(n_4458), .Z(n_4457));
   XOR2_X1 i_3948 (.A(n_1952), .B(n_4459), .Z(n_4458));
   XNOR2_X1 i_3949 (.A(n_1937), .B(n_4463), .ZN(n_4459));
   INV_X1 i_3950 (.A(n_4463), .ZN(n_4462));
   AOI21_X1 i_3951 (.A(n_1836), .B1(n_1835), .B2(n_4622), .ZN(n_4463));
   INV_X1 i_3952 (.A(n_4464), .ZN(n_1879));
   AOI21_X1 i_3953 (.A(n_1876), .B1(n_1875), .B2(n_4552), .ZN(n_4464));
   INV_X1 i_3954 (.A(n_4465), .ZN(n_1874));
   AOI21_X1 i_3955 (.A(n_1871), .B1(n_1870), .B2(n_4553), .ZN(n_4465));
   XNOR2_X1 i_3956 (.A(n_1967), .B(n_4467), .ZN(n_1969));
   INV_X1 i_3957 (.A(n_4467), .ZN(n_4466));
   AOI21_X1 i_3958 (.A(n_1861), .B1(n_1860), .B2(n_4558), .ZN(n_4467));
   INV_X1 i_3959 (.A(n_4469), .ZN(n_1869));
   AOI21_X1 i_3960 (.A(n_1866), .B1(n_1865), .B2(n_4568), .ZN(n_4469));
   XNOR2_X1 i_3961 (.A(n_1957), .B(n_4471), .ZN(n_1959));
   INV_X1 i_3962 (.A(n_4471), .ZN(n_4470));
   AOI21_X1 i_3963 (.A(n_1841), .B1(n_1840), .B2(n_4607), .ZN(n_4471));
   XOR2_X1 i_3964 (.A(n_1942), .B(n_4472), .Z(n_1944));
   XOR2_X1 i_3965 (.A(n_4475), .B(n_4473), .Z(n_4472));
   NAND2_X1 i_3966 (.A1(inputB[4]), .A2(inputA[15]), .ZN(n_4473));
   NAND2_X1 i_3967 (.A1(n_4478), .A2(n_4476), .ZN(n_4475));
   INV_X1 i_3968 (.A(n_4477), .ZN(n_4476));
   AOI22_X1 i_3969 (.A1(inputB[2]), .A2(inputA[17]), .B1(inputB[3]), .B2(
      inputA[16]), .ZN(n_4477));
   NAND2_X1 i_3970 (.A1(n_4611), .A2(n_4479), .ZN(n_4478));
   INV_X1 i_3971 (.A(n_4480), .ZN(n_4479));
   NAND2_X1 i_3972 (.A1(inputB[3]), .A2(inputA[17]), .ZN(n_4480));
   XOR2_X1 i_3973 (.A(n_1947), .B(n_4483), .Z(n_1949));
   XNOR2_X1 i_3974 (.A(n_4491), .B(n_4484), .ZN(n_4483));
   NOR2_X1 i_3975 (.A1(n_4490), .A2(n_4485), .ZN(n_4484));
   INV_X1 i_3976 (.A(n_4486), .ZN(n_4485));
   NAND3_X1 i_3977 (.A1(inputB[11]), .A2(inputA[7]), .A3(n_4487), .ZN(n_4486));
   INV_X1 i_3978 (.A(n_4488), .ZN(n_4487));
   NAND2_X1 i_3979 (.A1(inputB[12]), .A2(inputA[8]), .ZN(n_4488));
   AOI22_X1 i_3980 (.A1(inputB[11]), .A2(inputA[8]), .B1(inputB[12]), .B2(
      inputA[7]), .ZN(n_4490));
   NAND2_X1 i_3981 (.A1(inputB[13]), .A2(inputA[6]), .ZN(n_4491));
   INV_X1 i_3982 (.A(n_4492), .ZN(n_1859));
   AOI21_X1 i_3983 (.A(n_1856), .B1(n_1855), .B2(n_4600), .ZN(n_4492));
   INV_X1 i_3984 (.A(n_4493), .ZN(n_1854));
   AOI21_X1 i_3985 (.A(n_1851), .B1(n_1850), .B2(n_4602), .ZN(n_4493));
   INV_X1 i_3986 (.A(n_4494), .ZN(n_1849));
   AOI21_X1 i_3987 (.A(n_1846), .B1(n_1845), .B2(n_4573), .ZN(n_4494));
   XOR2_X1 i_3988 (.A(n_1932), .B(n_4496), .Z(n_1934));
   AOI21_X1 i_3989 (.A(n_4588), .B1(n_4587), .B2(n_4578), .ZN(n_4496));
   XOR2_X1 i_3990 (.A(n_4498), .B(n_4497), .Z(n_1884));
   NAND2_X1 i_3991 (.A1(inputB[19]), .A2(inputA[0]), .ZN(n_4497));
   NAND2_X1 i_3992 (.A1(n_4500), .A2(n_4499), .ZN(n_4498));
   NAND3_X1 i_3993 (.A1(inputB[17]), .A2(inputA[2]), .A3(n_4504), .ZN(n_4499));
   INV_X1 i_3994 (.A(n_4501), .ZN(n_4500));
   AOI21_X1 i_3995 (.A(n_4504), .B1(inputB[17]), .B2(inputA[2]), .ZN(n_4501));
   AND2_X1 i_3996 (.A1(inputB[18]), .A2(inputA[1]), .ZN(n_4504));
   XOR2_X1 i_3997 (.A(n_4506), .B(n_4505), .Z(n_1891));
   NAND2_X1 i_3998 (.A1(inputB[16]), .A2(inputA[3]), .ZN(n_4505));
   NAND2_X1 i_3999 (.A1(n_4508), .A2(n_4507), .ZN(n_4506));
   NAND3_X1 i_4000 (.A1(inputB[15]), .A2(inputA[5]), .A3(n_4635), .ZN(n_4507));
   INV_X1 i_4001 (.A(n_4509), .ZN(n_4508));
   AOI22_X1 i_4002 (.A1(inputB[14]), .A2(inputA[5]), .B1(inputB[15]), .B2(
      inputA[4]), .ZN(n_4509));
   XOR2_X1 i_4003 (.A(n_4511), .B(n_4510), .Z(n_1905));
   NAND2_X1 i_4004 (.A1(inputB[10]), .A2(inputA[9]), .ZN(n_4510));
   NAND2_X1 i_4005 (.A1(n_4513), .A2(n_4512), .ZN(n_4511));
   NAND3_X1 i_4006 (.A1(inputB[8]), .A2(inputA[11]), .A3(n_4517), .ZN(n_4512));
   INV_X1 i_4007 (.A(n_4514), .ZN(n_4513));
   AOI21_X1 i_4008 (.A(n_4517), .B1(inputB[8]), .B2(inputA[11]), .ZN(n_4514));
   AND2_X1 i_4009 (.A1(inputB[9]), .A2(inputA[10]), .ZN(n_4517));
   XOR2_X1 i_4010 (.A(n_4523), .B(n_4518), .Z(n_1912));
   NAND2_X1 i_4012 (.A1(inputB[7]), .A2(inputA[12]), .ZN(n_4518));
   NAND2_X1 i_4013 (.A1(n_4529), .A2(n_4528), .ZN(n_4523));
   NAND3_X1 i_4014 (.A1(inputB[6]), .A2(inputA[14]), .A3(n_4650), .ZN(n_4528));
   INV_X1 i_4016 (.A(n_4533), .ZN(n_4529));
   AOI22_X1 i_4017 (.A1(inputB[5]), .A2(inputA[14]), .B1(inputB[6]), .B2(
      inputA[13]), .ZN(n_4533));
   XOR2_X1 i_4018 (.A(n_4537), .B(n_4534), .Z(n_1925));
   AOI22_X1 i_4020 (.A1(n_4758), .A2(n_4612), .B1(n_4610), .B2(n_4608), .ZN(
      n_4534));
   AOI21_X1 i_4021 (.A(n_4538), .B1(n_4614), .B2(n_4543), .ZN(n_4537));
   AOI22_X1 i_4022 (.A1(inputB[1]), .A2(inputA[18]), .B1(inputB[0]), .B2(
      inputA[19]), .ZN(n_4538));
   AND2_X1 i_4024 (.A1(inputB[1]), .A2(inputA[19]), .ZN(n_4543));
   NAND2_X1 i_4025 (.A1(n_4616), .A2(n_4548), .ZN(n_1830));
   NAND2_X1 i_4026 (.A1(n_4617), .A2(n_4614), .ZN(n_4548));
   OAI21_X1 i_4028 (.A(n_4625), .B1(n_4629), .B2(n_4623), .ZN(n_1788));
   OAI21_X1 i_4029 (.A(n_4632), .B1(n_4634), .B2(n_4630), .ZN(n_1795));
   OAI21_X1 i_4030 (.A(n_4638), .B1(n_4642), .B2(n_4636), .ZN(n_1809));
   OAI21_X1 i_4032 (.A(n_4645), .B1(n_4649), .B2(n_4643), .ZN(n_1816));
   XOR2_X1 i_4033 (.A(n_1875), .B(n_4552), .Z(n_1877));
   XOR2_X1 i_4034 (.A(n_1870), .B(n_4553), .Z(n_4552));
   XNOR2_X1 i_4036 (.A(n_1860), .B(n_4559), .ZN(n_4553));
   INV_X1 i_4037 (.A(n_4559), .ZN(n_4558));
   AOI21_X1 i_4038 (.A(n_1764), .B1(n_1763), .B2(n_4694), .ZN(n_4559));
   INV_X1 i_4040 (.A(n_4562), .ZN(n_1782));
   AOI21_X1 i_4041 (.A(n_1779), .B1(n_1778), .B2(n_4563), .ZN(n_4562));
   XNOR2_X1 i_4042 (.A(n_1773), .B(n_4598), .ZN(n_4563));
   XOR2_X1 i_4044 (.A(n_1865), .B(n_4568), .Z(n_1867));
   XOR2_X1 i_4045 (.A(n_1845), .B(n_4573), .Z(n_4568));
   XNOR2_X1 i_4046 (.A(n_4583), .B(n_4578), .ZN(n_4573));
   NAND2_X1 i_4048 (.A1(inputB[12]), .A2(inputA[6]), .ZN(n_4578));
   NOR2_X1 i_4049 (.A1(n_4588), .A2(n_4584), .ZN(n_4583));
   INV_X1 i_4050 (.A(n_4587), .ZN(n_4584));
   NAND3_X1 i_4052 (.A1(inputB[11]), .A2(inputA[8]), .A3(n_4743), .ZN(n_4587));
   AOI22_X1 i_4053 (.A1(inputB[10]), .A2(inputA[8]), .B1(inputB[11]), .B2(
      inputA[7]), .ZN(n_4588));
   INV_X1 i_4054 (.A(n_4593), .ZN(n_1777));
   AOI21_X1 i_4056 (.A(n_1774), .B1(n_1773), .B2(n_4595), .ZN(n_4593));
   INV_X1 i_4057 (.A(n_4598), .ZN(n_4595));
   AOI21_X1 i_4058 (.A(n_1680), .B1(n_1679), .B2(n_4765), .ZN(n_4598));
   INV_X1 i_4060 (.A(n_4599), .ZN(n_1772));
   AOI21_X1 i_4061 (.A(n_1769), .B1(n_1768), .B2(n_4660), .ZN(n_4599));
   XNOR2_X1 i_4062 (.A(n_1855), .B(n_4601), .ZN(n_1857));
   INV_X1 i_4064 (.A(n_4601), .ZN(n_4600));
   AOI21_X1 i_4065 (.A(n_1754), .B1(n_1753), .B2(n_4705), .ZN(n_4601));
   XNOR2_X1 i_4066 (.A(n_1850), .B(n_4603), .ZN(n_1852));
   INV_X1 i_4068 (.A(n_4603), .ZN(n_4602));
   AOI21_X1 i_4069 (.A(n_1744), .B1(n_1743), .B2(n_4700), .ZN(n_4603));
   INV_X1 i_4070 (.A(n_4604), .ZN(n_1762));
   AOI21_X1 i_4072 (.A(n_1759), .B1(n_1758), .B2(n_4699), .ZN(n_4604));
   XOR2_X1 i_4073 (.A(n_1840), .B(n_4607), .Z(n_1842));
   XOR2_X1 i_4074 (.A(n_4609), .B(n_4608), .Z(n_4607));
   NAND2_X1 i_4076 (.A1(inputB[3]), .A2(inputA[15]), .ZN(n_4608));
   OAI21_X1 i_4077 (.A(n_4610), .B1(n_4755), .B2(n_4611), .ZN(n_4609));
   NAND2_X1 i_4078 (.A1(n_4755), .A2(n_4611), .ZN(n_4610));
   INV_X1 i_4079 (.A(n_4612), .ZN(n_4611));
   NAND2_X1 i_4080 (.A1(inputB[2]), .A2(inputA[16]), .ZN(n_4612));
   INV_X1 i_4081 (.A(n_4613), .ZN(n_1752));
   AOI21_X1 i_4082 (.A(n_1749), .B1(n_1748), .B2(n_4665), .ZN(n_4613));
   XOR2_X1 i_4083 (.A(n_4615), .B(n_4614), .Z(n_1829));
   AND2_X1 i_4084 (.A1(inputB[0]), .A2(inputA[18]), .ZN(n_4614));
   AND2_X1 i_4085 (.A1(n_4617), .A2(n_4616), .ZN(n_4615));
   NAND2_X1 i_4086 (.A1(n_4621), .A2(n_4618), .ZN(n_4616));
   OR2_X1 i_4087 (.A1(n_4621), .A2(n_4618), .ZN(n_4617));
   OAI21_X1 i_4088 (.A(n_4675), .B1(n_4680), .B2(n_4666), .ZN(n_4618));
   OAI21_X1 i_4089 (.A(n_4754), .B1(n_4760), .B2(n_4752), .ZN(n_4621));
   XOR2_X1 i_4090 (.A(n_1835), .B(n_4622), .Z(n_1837));
   OAI21_X1 i_4091 (.A(n_4715), .B1(n_4721), .B2(n_4709), .ZN(n_4622));
   XOR2_X1 i_4092 (.A(n_4624), .B(n_4623), .Z(n_1787));
   NAND2_X1 i_4093 (.A1(inputB[18]), .A2(inputA[0]), .ZN(n_4623));
   NAND2_X1 i_4094 (.A1(n_4628), .A2(n_4625), .ZN(n_4624));
   NAND4_X1 i_4095 (.A1(inputB[16]), .A2(inputA[2]), .A3(inputB[17]), .A4(
      inputA[1]), .ZN(n_4625));
   INV_X1 i_4096 (.A(n_4629), .ZN(n_4628));
   AOI22_X1 i_4097 (.A1(inputB[16]), .A2(inputA[2]), .B1(inputB[17]), .B2(
      inputA[1]), .ZN(n_4629));
   XOR2_X1 i_4098 (.A(n_4631), .B(n_4630), .Z(n_1794));
   NAND2_X1 i_4099 (.A1(inputB[15]), .A2(inputA[3]), .ZN(n_4630));
   NAND2_X1 i_4100 (.A1(n_4633), .A2(n_4632), .ZN(n_4631));
   NAND3_X1 i_4101 (.A1(inputB[13]), .A2(inputA[5]), .A3(n_4635), .ZN(n_4632));
   INV_X1 i_4102 (.A(n_4634), .ZN(n_4633));
   AOI21_X1 i_4103 (.A(n_4635), .B1(inputB[13]), .B2(inputA[5]), .ZN(n_4634));
   AND2_X1 i_4104 (.A1(inputB[14]), .A2(inputA[4]), .ZN(n_4635));
   XOR2_X1 i_4105 (.A(n_4637), .B(n_4636), .Z(n_1808));
   NAND2_X1 i_4106 (.A1(inputB[9]), .A2(inputA[9]), .ZN(n_4636));
   NAND2_X1 i_4107 (.A1(n_4639), .A2(n_4638), .ZN(n_4637));
   NAND4_X1 i_4108 (.A1(inputB[7]), .A2(inputA[11]), .A3(inputB[8]), .A4(
      inputA[10]), .ZN(n_4638));
   INV_X1 i_4109 (.A(n_4642), .ZN(n_4639));
   AOI22_X1 i_4110 (.A1(inputB[7]), .A2(inputA[11]), .B1(inputB[8]), .B2(
      inputA[10]), .ZN(n_4642));
   XOR2_X1 i_4111 (.A(n_4644), .B(n_4643), .Z(n_1815));
   NAND2_X1 i_4112 (.A1(inputB[6]), .A2(inputA[12]), .ZN(n_4643));
   NAND2_X1 i_4113 (.A1(n_4646), .A2(n_4645), .ZN(n_4644));
   NAND3_X1 i_4114 (.A1(inputB[4]), .A2(inputA[14]), .A3(n_4650), .ZN(n_4645));
   INV_X1 i_4115 (.A(n_4649), .ZN(n_4646));
   AOI21_X1 i_4116 (.A(n_4650), .B1(inputB[4]), .B2(inputA[14]), .ZN(n_4649));
   AND2_X1 i_4117 (.A1(inputB[5]), .A2(inputA[13]), .ZN(n_4650));
   INV_X1 i_4118 (.A(n_4651), .ZN(n_1742));
   AOI21_X1 i_4119 (.A(n_1739), .B1(n_1738), .B2(n_4730), .ZN(n_4651));
   OAI21_X1 i_4120 (.A(n_4737), .B1(n_4739), .B2(n_4735), .ZN(n_1699));
   AOI22_X1 i_4121 (.A1(n_4838), .A2(n_4744), .B1(n_4742), .B2(n_4740), .ZN(
      n_1713));
   OAI21_X1 i_4122 (.A(n_4747), .B1(n_4751), .B2(n_4745), .ZN(n_1720));
   INV_X1 i_4123 (.A(n_4654), .ZN(n_1693));
   AOI21_X1 i_4124 (.A(n_1690), .B1(n_1689), .B2(n_4655), .ZN(n_4654));
   XNOR2_X1 i_4125 (.A(n_1684), .B(n_4690), .ZN(n_4655));
   XOR2_X1 i_4126 (.A(n_1768), .B(n_4660), .Z(n_1770));
   XOR2_X1 i_4127 (.A(n_1748), .B(n_4665), .Z(n_4660));
   XOR2_X1 i_4128 (.A(n_4670), .B(n_4666), .Z(n_4665));
   NAND2_X1 i_4129 (.A1(inputB[5]), .A2(inputA[12]), .ZN(n_4666));
   NAND2_X1 i_4130 (.A1(n_4679), .A2(n_4675), .ZN(n_4670));
   NAND3_X1 i_4131 (.A1(inputB[4]), .A2(inputA[13]), .A3(n_4853), .ZN(n_4675));
   INV_X1 i_4132 (.A(n_4680), .ZN(n_4679));
   AOI21_X1 i_4133 (.A(n_4853), .B1(inputB[4]), .B2(inputA[13]), .ZN(n_4680));
   INV_X1 i_4134 (.A(n_4681), .ZN(n_1688));
   AOI21_X1 i_4135 (.A(n_1685), .B1(n_1684), .B2(n_4685), .ZN(n_4681));
   INV_X1 i_4136 (.A(n_4690), .ZN(n_4685));
   AOI21_X1 i_4137 (.A(n_1595), .B1(n_1594), .B2(n_4874), .ZN(n_4690));
   XNOR2_X1 i_4138 (.A(n_1763), .B(n_4695), .ZN(n_1765));
   INV_X1 i_4139 (.A(n_4695), .ZN(n_4694));
   AOI21_X1 i_4140 (.A(n_1665), .B1(n_1664), .B2(n_4779), .ZN(n_4695));
   XOR2_X1 i_4141 (.A(n_1758), .B(n_4699), .Z(n_1760));
   XNOR2_X1 i_4142 (.A(n_1743), .B(n_4701), .ZN(n_4699));
   INV_X1 i_4143 (.A(n_4701), .ZN(n_4700));
   AOI21_X1 i_4145 (.A(n_1655), .B1(n_1654), .B2(n_4807), .ZN(n_4701));
   XOR2_X1 i_4146 (.A(n_1753), .B(n_4705), .Z(n_1755));
   XOR2_X1 i_4147 (.A(n_4710), .B(n_4709), .Z(n_4705));
   NAND2_X1 i_4149 (.A1(inputB[14]), .A2(inputA[3]), .ZN(n_4709));
   NAND2_X1 i_4150 (.A1(n_4720), .A2(n_4715), .ZN(n_4710));
   NAND3_X1 i_4151 (.A1(inputB[13]), .A2(inputA[4]), .A3(n_4818), .ZN(n_4715));
   INV_X1 i_4153 (.A(n_4721), .ZN(n_4720));
   AOI21_X1 i_4154 (.A(n_4818), .B1(inputB[13]), .B2(inputA[4]), .ZN(n_4721));
   INV_X1 i_4155 (.A(n_4724), .ZN(n_1678));
   AOI21_X1 i_4157 (.A(n_1675), .B1(n_1674), .B2(n_4775), .ZN(n_4724));
   INV_X1 i_4158 (.A(n_4725), .ZN(n_1673));
   AOI21_X1 i_4159 (.A(n_1670), .B1(n_1669), .B2(n_4766), .ZN(n_4725));
   XOR2_X1 i_4161 (.A(n_1738), .B(n_4730), .Z(n_1740));
   OAI21_X1 i_4162 (.A(n_4833), .B1(n_4842), .B2(n_4828), .ZN(n_4730));
   INV_X1 i_4163 (.A(n_4732), .ZN(n_1663));
   AOI21_X1 i_4165 (.A(n_1660), .B1(n_1659), .B2(n_4789), .ZN(n_4732));
   XOR2_X1 i_4166 (.A(n_4736), .B(n_4735), .Z(n_1698));
   NAND2_X1 i_4167 (.A1(inputB[17]), .A2(inputA[0]), .ZN(n_4735));
   NAND2_X1 i_4169 (.A1(n_4738), .A2(n_4737), .ZN(n_4736));
   NAND3_X1 i_4170 (.A1(inputB[16]), .A2(inputA[1]), .A3(n_4772), .ZN(n_4737));
   INV_X1 i_4171 (.A(n_4739), .ZN(n_4738));
   AOI21_X1 i_4173 (.A(n_4772), .B1(inputB[16]), .B2(inputA[1]), .ZN(n_4739));
   XOR2_X1 i_4174 (.A(n_4741), .B(n_4740), .Z(n_1712));
   NAND2_X1 i_4175 (.A1(inputB[11]), .A2(inputA[6]), .ZN(n_4740));
   OAI21_X1 i_4177 (.A(n_4742), .B1(n_4834), .B2(n_4743), .ZN(n_4741));
   NAND2_X1 i_4178 (.A1(n_4834), .A2(n_4743), .ZN(n_4742));
   INV_X1 i_4179 (.A(n_4744), .ZN(n_4743));
   NAND2_X1 i_4181 (.A1(inputB[10]), .A2(inputA[7]), .ZN(n_4744));
   XOR2_X1 i_4182 (.A(n_4746), .B(n_4745), .Z(n_1719));
   NAND2_X1 i_4183 (.A1(inputB[8]), .A2(inputA[9]), .ZN(n_4745));
   NAND2_X1 i_4185 (.A1(n_4748), .A2(n_4747), .ZN(n_4746));
   NAND3_X1 i_4186 (.A1(inputB[7]), .A2(inputA[10]), .A3(n_4785), .ZN(n_4747));
   INV_X1 i_4187 (.A(n_4751), .ZN(n_4748));
   AOI21_X1 i_4189 (.A(n_4785), .B1(inputB[7]), .B2(inputA[10]), .ZN(n_4751));
   XOR2_X1 i_4190 (.A(n_4753), .B(n_4752), .Z(n_1733));
   NAND2_X1 i_4191 (.A1(inputB[2]), .A2(inputA[15]), .ZN(n_4752));
   NAND2_X1 i_4193 (.A1(n_4759), .A2(n_4754), .ZN(n_4753));
   NAND2_X1 i_4194 (.A1(n_4870), .A2(n_4755), .ZN(n_4754));
   INV_X1 i_4195 (.A(n_4758), .ZN(n_4755));
   NAND2_X1 i_4197 (.A1(inputB[1]), .A2(inputA[17]), .ZN(n_4758));
   INV_X1 i_4198 (.A(n_4760), .ZN(n_4759));
   AOI22_X1 i_4199 (.A1(inputB[0]), .A2(inputA[17]), .B1(inputB[1]), .B2(
      inputA[16]), .ZN(n_4760));
   OAI21_X1 i_4201 (.A(n_4865), .B1(n_4868), .B2(n_4858), .ZN(n_1648));
   OAI21_X1 i_4202 (.A(n_4769), .B1(n_4774), .B2(n_4767), .ZN(n_1614));
   OAI21_X1 i_4203 (.A(n_4817), .B1(n_4823), .B2(n_4808), .ZN(n_1621));
   OAI21_X1 i_4205 (.A(n_4784), .B1(n_4783), .B2(n_4780), .ZN(n_1635));
   OAI21_X1 i_4206 (.A(n_4849), .B1(n_4857), .B2(n_4843), .ZN(n_1642));
   INV_X1 i_4207 (.A(n_4761), .ZN(n_1608));
   AOI21_X1 i_4208 (.A(n_1605), .B1(n_1604), .B2(n_4762), .ZN(n_4761));
   XOR2_X1 i_4209 (.A(n_1599), .B(n_4764), .Z(n_4762));
   INV_X1 i_4210 (.A(n_4763), .ZN(n_1603));
   AOI21_X1 i_4211 (.A(n_1600), .B1(n_1599), .B2(n_4764), .ZN(n_4763));
   XOR2_X1 i_4212 (.A(n_1589), .B(n_4787), .Z(n_4764));
   XOR2_X1 i_4213 (.A(n_1679), .B(n_4765), .Z(n_1681));
   XOR2_X1 i_4214 (.A(n_1669), .B(n_4766), .Z(n_4765));
   XOR2_X1 i_4215 (.A(n_4768), .B(n_4767), .Z(n_4766));
   NAND2_X1 i_4216 (.A1(inputB[16]), .A2(inputA[0]), .ZN(n_4767));
   NAND2_X1 i_4217 (.A1(n_4773), .A2(n_4769), .ZN(n_4768));
   NAND3_X1 i_4218 (.A1(inputB[14]), .A2(inputA[1]), .A3(n_4772), .ZN(n_4769));
   AND2_X1 i_4219 (.A1(inputB[15]), .A2(inputA[2]), .ZN(n_4772));
   INV_X1 i_4220 (.A(n_4774), .ZN(n_4773));
   AOI22_X1 i_4221 (.A1(inputB[14]), .A2(inputA[2]), .B1(inputB[15]), .B2(
      inputA[1]), .ZN(n_4774));
   XNOR2_X1 i_4222 (.A(n_1674), .B(n_4776), .ZN(n_1676));
   INV_X1 i_4223 (.A(n_4776), .ZN(n_4775));
   AOI21_X1 i_4224 (.A(n_1580), .B1(n_1579), .B2(n_4886), .ZN(n_4776));
   XOR2_X1 i_4225 (.A(n_1664), .B(n_4779), .Z(n_1666));
   XOR2_X1 i_4226 (.A(n_4781), .B(n_4780), .Z(n_4779));
   NAND2_X1 i_4227 (.A1(inputB[7]), .A2(inputA[9]), .ZN(n_4780));
   NAND2_X1 i_4228 (.A1(n_4784), .A2(n_4782), .ZN(n_4781));
   INV_X1 i_4229 (.A(n_4783), .ZN(n_4782));
   AOI22_X1 i_4230 (.A1(inputB[5]), .A2(inputA[11]), .B1(inputB[6]), .B2(
      inputA[10]), .ZN(n_4783));
   NAND2_X1 i_4231 (.A1(n_4894), .A2(n_4785), .ZN(n_4784));
   AND2_X1 i_4232 (.A1(inputB[6]), .A2(inputA[11]), .ZN(n_4785));
   INV_X1 i_4233 (.A(n_4786), .ZN(n_1593));
   AOI21_X1 i_4234 (.A(n_1590), .B1(n_1589), .B2(n_4787), .ZN(n_4786));
   XOR2_X1 i_4235 (.A(n_4793), .B(n_4788), .Z(n_4787));
   OAI21_X1 i_4236 (.A(n_4794), .B1(n_4803), .B2(n_4802), .ZN(n_4788));
   XOR2_X1 i_4237 (.A(n_1659), .B(n_4789), .Z(n_1661));
   OAI21_X1 i_4238 (.A(n_4794), .B1(n_4798), .B2(n_4793), .ZN(n_4789));
   NAND2_X1 i_4239 (.A1(inputB[0]), .A2(inputA[15]), .ZN(n_4793));
   NAND2_X1 i_4240 (.A1(n_4803), .A2(n_4802), .ZN(n_4794));
   NOR2_X1 i_4241 (.A1(n_4803), .A2(n_4802), .ZN(n_4798));
   AOI21_X1 i_4242 (.A(n_5007), .B1(n_5006), .B2(n_5002), .ZN(n_4802));
   AOI21_X1 i_4243 (.A(n_5013), .B1(n_5014), .B2(n_5008), .ZN(n_4803));
   INV_X1 i_4244 (.A(n_4804), .ZN(n_1588));
   AOI21_X1 i_4245 (.A(n_1585), .B1(n_1584), .B2(n_4877), .ZN(n_4804));
   XOR2_X1 i_4246 (.A(n_1654), .B(n_4807), .Z(n_1656));
   OAI21_X1 i_4247 (.A(n_4906), .B1(n_4908), .B2(n_4904), .ZN(n_4807));
   XOR2_X1 i_4248 (.A(n_4813), .B(n_4808), .Z(n_1620));
   NAND2_X1 i_4249 (.A1(inputB[13]), .A2(inputA[3]), .ZN(n_4808));
   NAND2_X1 i_4250 (.A1(n_4819), .A2(n_4817), .ZN(n_4813));
   NAND2_X1 i_4251 (.A1(n_4909), .A2(n_4818), .ZN(n_4817));
   AND2_X1 i_4252 (.A1(inputB[12]), .A2(inputA[5]), .ZN(n_4818));
   INV_X1 i_4253 (.A(n_4823), .ZN(n_4819));
   AOI22_X1 i_4254 (.A1(inputB[11]), .A2(inputA[5]), .B1(inputB[12]), .B2(
      inputA[4]), .ZN(n_4823));
   XOR2_X1 i_4255 (.A(n_4832), .B(n_4828), .Z(n_1627));
   NAND2_X1 i_4256 (.A1(inputB[10]), .A2(inputA[6]), .ZN(n_4828));
   NAND2_X1 i_4257 (.A1(n_4839), .A2(n_4833), .ZN(n_4832));
   NAND2_X1 i_4258 (.A1(n_4915), .A2(n_4834), .ZN(n_4833));
   INV_X1 i_4259 (.A(n_4838), .ZN(n_4834));
   NAND2_X1 i_4260 (.A1(inputB[9]), .A2(inputA[8]), .ZN(n_4838));
   INV_X1 i_4261 (.A(n_4842), .ZN(n_4839));
   AOI22_X1 i_4262 (.A1(inputB[8]), .A2(inputA[8]), .B1(inputB[9]), .B2(
      inputA[7]), .ZN(n_4842));
   XOR2_X1 i_4263 (.A(n_4848), .B(n_4843), .Z(n_1641));
   NAND2_X1 i_4264 (.A1(inputB[4]), .A2(inputA[12]), .ZN(n_4843));
   NAND2_X1 i_4266 (.A1(n_4854), .A2(n_4849), .ZN(n_4848));
   NAND2_X1 i_4267 (.A1(n_4922), .A2(n_4853), .ZN(n_4849));
   AND2_X1 i_4268 (.A1(inputB[3]), .A2(inputA[14]), .ZN(n_4853));
   INV_X1 i_4270 (.A(n_4857), .ZN(n_4854));
   AOI22_X1 i_4271 (.A1(inputB[2]), .A2(inputA[14]), .B1(inputB[3]), .B2(
      inputA[13]), .ZN(n_4857));
   XOR2_X1 i_4272 (.A(n_4863), .B(n_4858), .Z(n_1647));
   NAND2_X1 i_4274 (.A1(inputB[1]), .A2(inputA[15]), .ZN(n_4858));
   OAI21_X1 i_4275 (.A(n_4865), .B1(n_4870), .B2(n_4869), .ZN(n_4863));
   NAND2_X1 i_4276 (.A1(n_4870), .A2(n_4869), .ZN(n_4865));
   NOR2_X1 i_4278 (.A1(n_4870), .A2(n_4869), .ZN(n_4868));
   AOI22_X1 i_4279 (.A1(n_5016), .A2(n_4926), .B1(n_4921), .B2(n_4919), .ZN(
      n_4869));
   AND2_X1 i_4280 (.A1(inputB[0]), .A2(inputA[16]), .ZN(n_4870));
   INV_X1 i_4282 (.A(n_4871), .ZN(n_1578));
   AOI21_X1 i_4283 (.A(n_1575), .B1(n_1574), .B2(n_4901), .ZN(n_4871));
   OAI21_X1 i_4284 (.A(n_4880), .B1(n_4882), .B2(n_4881), .ZN(n_1534));
   AOI22_X1 i_4286 (.A1(n_4941), .A2(n_4916), .B1(n_4914), .B2(n_4912), .ZN(
      n_1548));
   OAI21_X1 i_4287 (.A(n_4891), .B1(n_4893), .B2(n_4887), .ZN(n_1555));
   INV_X1 i_4288 (.A(n_4872), .ZN(n_1528));
   AOI21_X1 i_4290 (.A(n_1525), .B1(n_1524), .B2(n_4873), .ZN(n_4872));
   XOR2_X1 i_4291 (.A(n_1519), .B(n_4884), .Z(n_4873));
   XOR2_X1 i_4292 (.A(n_1594), .B(n_4874), .Z(n_1596));
   XOR2_X1 i_4294 (.A(n_1584), .B(n_4877), .Z(n_4874));
   XNOR2_X1 i_4295 (.A(n_4882), .B(n_4878), .ZN(n_4877));
   NOR2_X1 i_4296 (.A1(n_4881), .A2(n_4879), .ZN(n_4878));
   INV_X1 i_4298 (.A(n_4880), .ZN(n_4879));
   NAND3_X1 i_4299 (.A1(inputB[14]), .A2(inputA[2]), .A3(n_4994), .ZN(n_4880));
   AOI22_X1 i_4300 (.A1(inputB[13]), .A2(inputA[2]), .B1(inputB[14]), .B2(
      inputA[1]), .ZN(n_4881));
   NAND2_X1 i_4302 (.A1(inputB[15]), .A2(inputA[0]), .ZN(n_4882));
   INV_X1 i_4303 (.A(n_4883), .ZN(n_1523));
   AOI21_X1 i_4304 (.A(n_1520), .B1(n_1519), .B2(n_4884), .ZN(n_4883));
   XOR2_X1 i_4306 (.A(n_1504), .B(n_4899), .Z(n_4884));
   INV_X1 i_4307 (.A(n_4885), .ZN(n_1518));
   AOI21_X1 i_4308 (.A(n_1515), .B1(n_1514), .B2(n_4961), .ZN(n_4885));
   XOR2_X1 i_4310 (.A(n_1579), .B(n_4886), .Z(n_1581));
   XOR2_X1 i_4311 (.A(n_4888), .B(n_4887), .Z(n_4886));
   NAND2_X1 i_4312 (.A1(inputB[6]), .A2(inputA[9]), .ZN(n_4887));
   NAND2_X1 i_4314 (.A1(n_4892), .A2(n_4891), .ZN(n_4888));
   NAND3_X1 i_4315 (.A1(inputB[4]), .A2(inputA[11]), .A3(n_4894), .ZN(n_4891));
   INV_X1 i_4316 (.A(n_4893), .ZN(n_4892));
   AOI21_X1 i_4318 (.A(n_4894), .B1(inputB[4]), .B2(inputA[11]), .ZN(n_4893));
   AND2_X1 i_4319 (.A1(inputB[5]), .A2(inputA[10]), .ZN(n_4894));
   INV_X1 i_4320 (.A(n_4895), .ZN(n_1513));
   AOI21_X1 i_4322 (.A(n_1510), .B1(n_1509), .B2(n_4967), .ZN(n_4895));
   INV_X1 i_4323 (.A(n_4898), .ZN(n_1508));
   AOI21_X1 i_4324 (.A(n_1505), .B1(n_1504), .B2(n_4899), .ZN(n_4898));
   XNOR2_X1 i_4326 (.A(n_4932), .B(n_4900), .ZN(n_4899));
   AOI21_X1 i_4327 (.A(n_4942), .B1(n_5096), .B2(n_4936), .ZN(n_4900));
   XOR2_X1 i_4328 (.A(n_1574), .B(n_4901), .Z(n_1576));
   NAND2_X1 i_4329 (.A1(n_4993), .A2(n_4902), .ZN(n_4901));
   NAND2_X1 i_4330 (.A1(n_4991), .A2(n_4985), .ZN(n_4902));
   INV_X1 i_4331 (.A(n_4903), .ZN(n_1503));
   AOI21_X1 i_4332 (.A(n_1500), .B1(n_1499), .B2(n_4962), .ZN(n_4903));
   XOR2_X1 i_4333 (.A(n_4905), .B(n_4904), .Z(n_1540));
   NAND2_X1 i_4334 (.A1(inputB[12]), .A2(inputA[3]), .ZN(n_4904));
   NAND2_X1 i_4335 (.A1(n_4907), .A2(n_4906), .ZN(n_4905));
   NAND3_X1 i_4336 (.A1(inputB[10]), .A2(inputA[5]), .A3(n_4909), .ZN(n_4906));
   INV_X1 i_4337 (.A(n_4908), .ZN(n_4907));
   AOI21_X1 i_4338 (.A(n_4909), .B1(inputB[10]), .B2(inputA[5]), .ZN(n_4908));
   AND2_X1 i_4339 (.A1(inputB[11]), .A2(inputA[4]), .ZN(n_4909));
   XOR2_X1 i_4340 (.A(n_4913), .B(n_4912), .Z(n_1547));
   NAND2_X1 i_4341 (.A1(inputB[9]), .A2(inputA[6]), .ZN(n_4912));
   OAI21_X1 i_4342 (.A(n_4914), .B1(n_4936), .B2(n_4915), .ZN(n_4913));
   NAND2_X1 i_4343 (.A1(n_4936), .A2(n_4915), .ZN(n_4914));
   INV_X1 i_4344 (.A(n_4916), .ZN(n_4915));
   NAND2_X1 i_4345 (.A1(inputB[8]), .A2(inputA[7]), .ZN(n_4916));
   XOR2_X1 i_4346 (.A(n_4920), .B(n_4919), .Z(n_1561));
   NAND2_X1 i_4347 (.A1(inputB[3]), .A2(inputA[12]), .ZN(n_4919));
   OAI21_X1 i_4348 (.A(n_4921), .B1(n_5015), .B2(n_4922), .ZN(n_4920));
   NAND2_X1 i_4349 (.A1(n_5015), .A2(n_4922), .ZN(n_4921));
   INV_X1 i_4350 (.A(n_4926), .ZN(n_4922));
   NAND2_X1 i_4351 (.A1(inputB[2]), .A2(inputA[13]), .ZN(n_4926));
   INV_X1 i_4352 (.A(n_4931), .ZN(n_1498));
   AOI21_X1 i_4353 (.A(n_1495), .B1(n_1494), .B2(n_4971), .ZN(n_4931));
   OAI21_X1 i_4354 (.A(n_4999), .B1(n_5001), .B2(n_4997), .ZN(n_1469));
   OAI21_X1 i_4355 (.A(n_4935), .B1(n_4942), .B2(n_4932), .ZN(n_1476));
   NAND2_X1 i_4356 (.A1(inputB[8]), .A2(inputA[6]), .ZN(n_4932));
   NAND2_X1 i_4357 (.A1(n_5096), .A2(n_4936), .ZN(n_4935));
   INV_X1 i_4358 (.A(n_4941), .ZN(n_4936));
   NAND2_X1 i_4359 (.A1(inputB[7]), .A2(inputA[8]), .ZN(n_4941));
   AOI22_X1 i_4360 (.A1(inputB[6]), .A2(inputA[8]), .B1(inputB[7]), .B2(
      inputA[7]), .ZN(n_4942));
   INV_X1 i_4361 (.A(n_4946), .ZN(n_1456));
   AOI21_X1 i_4362 (.A(n_1453), .B1(n_1452), .B2(n_4950), .ZN(n_4946));
   INV_X1 i_4363 (.A(n_4951), .ZN(n_4950));
   AOI21_X1 i_4364 (.A(n_1385), .B1(n_1384), .B2(n_4956), .ZN(n_4951));
   XOR2_X1 i_4365 (.A(n_1379), .B(n_5029), .Z(n_4956));
   INV_X1 i_4366 (.A(n_4957), .ZN(n_1451));
   AOI21_X1 i_4367 (.A(n_1448), .B1(n_1447), .B2(n_5019), .ZN(n_4957));
   XOR2_X1 i_4368 (.A(n_1514), .B(n_4961), .Z(n_1516));
   XNOR2_X1 i_4369 (.A(n_1499), .B(n_4966), .ZN(n_4961));
   INV_X1 i_4370 (.A(n_4966), .ZN(n_4962));
   AOI22_X1 i_4371 (.A1(n_5105), .A2(n_5102), .B1(n_5101), .B2(n_5097), .ZN(
      n_4966));
   XOR2_X1 i_4372 (.A(n_1509), .B(n_4967), .Z(n_1511));
   XOR2_X1 i_4373 (.A(n_1494), .B(n_4971), .Z(n_4967));
   OAI21_X1 i_4374 (.A(n_5067), .B1(n_5076), .B2(n_5061), .ZN(n_4971));
   INV_X1 i_4375 (.A(n_4976), .ZN(n_1446));
   AOI21_X1 i_4376 (.A(n_1443), .B1(n_1442), .B2(n_5030), .ZN(n_4976));
   INV_X1 i_4377 (.A(n_4977), .ZN(n_1436));
   AOI21_X1 i_4378 (.A(n_1433), .B1(n_1432), .B2(n_5020), .ZN(n_4977));
   INV_X1 i_4379 (.A(n_4981), .ZN(n_1441));
   AOI21_X1 i_4380 (.A(n_1438), .B1(n_1437), .B2(n_5036), .ZN(n_4981));
   XOR2_X1 i_4381 (.A(n_4986), .B(n_4985), .Z(n_1461));
   AND2_X1 i_4382 (.A1(inputB[14]), .A2(inputA[0]), .ZN(n_4985));
   AND2_X1 i_4383 (.A1(n_4993), .A2(n_4991), .ZN(n_4986));
   NAND2_X1 i_4384 (.A1(n_5047), .A2(n_4996), .ZN(n_4991));
   NAND2_X1 i_4385 (.A1(n_5046), .A2(n_4994), .ZN(n_4993));
   INV_X1 i_4386 (.A(n_4996), .ZN(n_4994));
   NAND2_X1 i_4388 (.A1(inputB[13]), .A2(inputA[1]), .ZN(n_4996));
   XOR2_X1 i_4389 (.A(n_4998), .B(n_4997), .Z(n_1468));
   NAND2_X1 i_4390 (.A1(inputB[11]), .A2(inputA[3]), .ZN(n_4997));
   NAND2_X1 i_4392 (.A1(n_5000), .A2(n_4999), .ZN(n_4998));
   NAND4_X1 i_4393 (.A1(inputB[9]), .A2(inputA[5]), .A3(inputB[10]), .A4(
      inputA[4]), .ZN(n_4999));
   INV_X1 i_4394 (.A(n_5001), .ZN(n_5000));
   AOI22_X1 i_4396 (.A1(inputB[9]), .A2(inputA[5]), .B1(inputB[10]), .B2(
      inputA[4]), .ZN(n_5001));
   XNOR2_X1 i_4397 (.A(n_5004), .B(n_5002), .ZN(n_1482));
   NAND2_X1 i_4398 (.A1(inputB[5]), .A2(inputA[9]), .ZN(n_5002));
   NOR2_X1 i_4400 (.A1(n_5007), .A2(n_5005), .ZN(n_5004));
   INV_X1 i_4401 (.A(n_5006), .ZN(n_5005));
   NAND3_X1 i_4402 (.A1(inputB[4]), .A2(inputA[10]), .A3(n_5027), .ZN(n_5006));
   AOI21_X1 i_4404 (.A(n_5027), .B1(inputB[4]), .B2(inputA[10]), .ZN(n_5007));
   XOR2_X1 i_4405 (.A(n_5009), .B(n_5008), .Z(n_1489));
   NAND2_X1 i_4406 (.A1(inputB[2]), .A2(inputA[12]), .ZN(n_5008));
   NAND2_X1 i_4408 (.A1(n_5014), .A2(n_5012), .ZN(n_5009));
   INV_X1 i_4409 (.A(n_5013), .ZN(n_5012));
   AOI22_X1 i_4410 (.A1(inputB[1]), .A2(inputA[13]), .B1(inputB[0]), .B2(
      inputA[14]), .ZN(n_5013));
   NAND2_X1 i_4412 (.A1(n_5105), .A2(n_5015), .ZN(n_5014));
   INV_X1 i_4413 (.A(n_5016), .ZN(n_5015));
   NAND2_X1 i_4414 (.A1(inputB[1]), .A2(inputA[14]), .ZN(n_5016));
   INV_X1 i_4416 (.A(n_5017), .ZN(n_1431));
   AOI21_X1 i_4417 (.A(n_1428), .B1(n_1427), .B2(n_5051), .ZN(n_5017));
   OAI21_X1 i_4418 (.A(n_5042), .B1(n_5041), .B2(n_5037), .ZN(n_1394));
   OAI21_X1 i_4420 (.A(n_5086), .B1(n_5095), .B2(n_5081), .ZN(n_1408));
   OAI21_X1 i_4421 (.A(n_5026), .B1(n_5025), .B2(n_5021), .ZN(n_1415));
   XOR2_X1 i_4422 (.A(n_1447), .B(n_5019), .Z(n_1449));
   XOR2_X1 i_4424 (.A(n_1432), .B(n_5020), .Z(n_5019));
   XOR2_X1 i_4425 (.A(n_5022), .B(n_5021), .Z(n_5020));
   NAND2_X1 i_4426 (.A1(inputB[4]), .A2(inputA[9]), .ZN(n_5021));
   NAND2_X1 i_4428 (.A1(n_5026), .A2(n_5023), .ZN(n_5022));
   INV_X1 i_4429 (.A(n_5025), .ZN(n_5023));
   AOI22_X1 i_4430 (.A1(inputB[2]), .A2(inputA[11]), .B1(inputB[3]), .B2(
      inputA[10]), .ZN(n_5025));
   NAND3_X1 i_4432 (.A1(inputB[2]), .A2(inputA[10]), .A3(n_5027), .ZN(n_5026));
   AND2_X1 i_4433 (.A1(inputB[3]), .A2(inputA[11]), .ZN(n_5027));
   INV_X1 i_4434 (.A(n_5028), .ZN(n_1383));
   AOI21_X1 i_4436 (.A(n_1380), .B1(n_1379), .B2(n_5029), .ZN(n_5028));
   XOR2_X1 i_4437 (.A(n_1369), .B(n_5034), .Z(n_5029));
   XNOR2_X1 i_4438 (.A(n_1442), .B(n_5033), .ZN(n_1444));
   INV_X1 i_4440 (.A(n_5033), .ZN(n_5030));
   AOI21_X1 i_4441 (.A(n_1370), .B1(n_1369), .B2(n_5034), .ZN(n_5033));
   XNOR2_X1 i_4442 (.A(n_5111), .B(n_5035), .ZN(n_5034));
   AOI21_X1 i_4444 (.A(n_5116), .B1(n_5229), .B2(n_5115), .ZN(n_5035));
   XOR2_X1 i_4445 (.A(n_1437), .B(n_5036), .Z(n_1439));
   XOR2_X1 i_4446 (.A(n_5038), .B(n_5037), .Z(n_5036));
   NAND2_X1 i_4447 (.A1(inputB[13]), .A2(inputA[0]), .ZN(n_5037));
   NAND2_X1 i_4448 (.A1(n_5042), .A2(n_5040), .ZN(n_5038));
   INV_X1 i_4449 (.A(n_5041), .ZN(n_5040));
   AOI22_X1 i_4450 (.A1(inputB[11]), .A2(inputA[2]), .B1(inputB[12]), .B2(
      inputA[1]), .ZN(n_5041));
   NAND2_X1 i_4451 (.A1(n_5142), .A2(n_5046), .ZN(n_5042));
   INV_X1 i_4452 (.A(n_5047), .ZN(n_5046));
   NAND2_X1 i_4453 (.A1(inputB[12]), .A2(inputA[2]), .ZN(n_5047));
   INV_X1 i_4454 (.A(n_5050), .ZN(n_1378));
   AOI21_X1 i_4455 (.A(n_1375), .B1(n_1374), .B2(n_5119), .ZN(n_5050));
   XOR2_X1 i_4456 (.A(n_1427), .B(n_5051), .Z(n_1429));
   OAI21_X1 i_4457 (.A(n_5139), .B1(n_5141), .B2(n_5136), .ZN(n_5051));
   INV_X1 i_4458 (.A(n_5056), .ZN(n_1368));
   AOI21_X1 i_4459 (.A(n_1365), .B1(n_1364), .B2(n_5134), .ZN(n_5056));
   XOR2_X1 i_4460 (.A(n_5066), .B(n_5061), .Z(n_1400));
   NAND2_X1 i_4461 (.A1(inputB[10]), .A2(inputA[3]), .ZN(n_5061));
   NAND2_X1 i_4462 (.A1(n_5071), .A2(n_5067), .ZN(n_5066));
   NAND3_X1 i_4463 (.A1(inputB[9]), .A2(inputA[4]), .A3(n_5115), .ZN(n_5067));
   INV_X1 i_4464 (.A(n_5076), .ZN(n_5071));
   AOI21_X1 i_4465 (.A(n_5115), .B1(inputB[9]), .B2(inputA[4]), .ZN(n_5076));
   XOR2_X1 i_4466 (.A(n_5082), .B(n_5081), .Z(n_1407));
   NAND2_X1 i_4467 (.A1(inputB[7]), .A2(inputA[6]), .ZN(n_5081));
   NAND2_X1 i_4468 (.A1(n_5091), .A2(n_5086), .ZN(n_5082));
   NAND3_X1 i_4469 (.A1(inputB[5]), .A2(inputA[8]), .A3(n_5096), .ZN(n_5086));
   INV_X1 i_4470 (.A(n_5095), .ZN(n_5091));
   AOI21_X1 i_4471 (.A(n_5096), .B1(inputB[5]), .B2(inputA[8]), .ZN(n_5095));
   AND2_X1 i_4472 (.A1(inputB[6]), .A2(inputA[7]), .ZN(n_5096));
   XOR2_X1 i_4473 (.A(n_5101), .B(n_5097), .Z(n_1420));
   OAI22_X1 i_4474 (.A1(n_5234), .A2(n_5155), .B1(n_5153), .B2(n_5149), .ZN(
      n_5097));
   XNOR2_X1 i_4475 (.A(n_5106), .B(n_5102), .ZN(n_5101));
   AND2_X1 i_4476 (.A1(inputB[1]), .A2(inputA[12]), .ZN(n_5102));
   INV_X1 i_4477 (.A(n_5106), .ZN(n_5105));
   NAND2_X1 i_4478 (.A1(inputB[0]), .A2(inputA[13]), .ZN(n_5106));
   OAI21_X1 i_4479 (.A(n_5122), .B1(n_5123), .B2(n_5120), .ZN(n_1359));
   OAI21_X1 i_4480 (.A(n_5113), .B1(n_5116), .B2(n_5111), .ZN(n_1338));
   NAND2_X1 i_4481 (.A1(inputB[9]), .A2(inputA[3]), .ZN(n_5111));
   NAND2_X1 i_4482 (.A1(n_5229), .A2(n_5115), .ZN(n_5113));
   AND2_X1 i_4483 (.A1(inputB[8]), .A2(inputA[5]), .ZN(n_5115));
   AOI22_X1 i_4484 (.A1(inputB[7]), .A2(inputA[5]), .B1(inputB[8]), .B2(
      inputA[4]), .ZN(n_5116));
   OAI21_X1 i_4485 (.A(n_5146), .B1(n_5148), .B2(n_5143), .ZN(n_1345));
   INV_X1 i_4486 (.A(n_5117), .ZN(n_1325));
   AOI21_X1 i_4487 (.A(n_1322), .B1(n_1321), .B2(n_5118), .ZN(n_5117));
   XNOR2_X1 i_4488 (.A(n_1316), .B(n_5129), .ZN(n_5118));
   XOR2_X1 i_4489 (.A(n_1374), .B(n_5119), .Z(n_1376));
   XOR2_X1 i_4490 (.A(n_5121), .B(n_5120), .Z(n_5119));
   NAND2_X1 i_4491 (.A1(inputB[0]), .A2(inputA[12]), .ZN(n_5120));
   OAI21_X1 i_4492 (.A(n_5122), .B1(n_5126), .B2(n_5125), .ZN(n_5121));
   NAND2_X1 i_4493 (.A1(n_5126), .A2(n_5125), .ZN(n_5122));
   NOR2_X1 i_4494 (.A1(n_5126), .A2(n_5125), .ZN(n_5123));
   OAI22_X1 i_4495 (.A1(n_5279), .A2(n_5234), .B1(n_5236), .B2(n_5232), .ZN(
      n_5125));
   OAI21_X1 i_4496 (.A(n_5177), .B1(n_5172), .B2(n_5163), .ZN(n_5126));
   INV_X1 i_4497 (.A(n_5127), .ZN(n_1320));
   AOI21_X1 i_4498 (.A(n_1317), .B1(n_1316), .B2(n_5128), .ZN(n_5127));
   INV_X1 i_4499 (.A(n_5129), .ZN(n_5128));
   AOI21_X1 i_4500 (.A(n_1262), .B1(n_1261), .B2(n_5160), .ZN(n_5129));
   INV_X1 i_4501 (.A(n_5132), .ZN(n_1315));
   AOI21_X1 i_4502 (.A(n_1312), .B1(n_1311), .B2(n_5182), .ZN(n_5132));
   INV_X1 i_4503 (.A(n_5133), .ZN(n_1310));
   AOI21_X1 i_4504 (.A(n_1307), .B1(n_1306), .B2(n_5162), .ZN(n_5133));
   XNOR2_X1 i_4506 (.A(n_1364), .B(n_5135), .ZN(n_1366));
   INV_X1 i_4507 (.A(n_5135), .ZN(n_5134));
   AOI21_X1 i_4508 (.A(n_1302), .B1(n_1301), .B2(n_5196), .ZN(n_5135));
   XOR2_X1 i_4510 (.A(n_5138), .B(n_5136), .Z(n_1330));
   NAND2_X1 i_4511 (.A1(inputB[12]), .A2(inputA[0]), .ZN(n_5136));
   NAND2_X1 i_4512 (.A1(n_5140), .A2(n_5139), .ZN(n_5138));
   NAND3_X1 i_4514 (.A1(inputB[10]), .A2(inputA[2]), .A3(n_5142), .ZN(n_5139));
   INV_X1 i_4515 (.A(n_5141), .ZN(n_5140));
   AOI21_X1 i_4516 (.A(n_5142), .B1(inputB[10]), .B2(inputA[2]), .ZN(n_5141));
   AND2_X1 i_4518 (.A1(inputB[11]), .A2(inputA[1]), .ZN(n_5142));
   XOR2_X1 i_4519 (.A(n_5144), .B(n_5143), .Z(n_1344));
   NAND2_X1 i_4520 (.A1(inputB[6]), .A2(inputA[6]), .ZN(n_5143));
   NAND2_X1 i_4522 (.A1(n_5147), .A2(n_5146), .ZN(n_5144));
   NAND3_X1 i_4523 (.A1(inputB[5]), .A2(inputA[7]), .A3(n_5181), .ZN(n_5146));
   INV_X1 i_4524 (.A(n_5148), .ZN(n_5147));
   AOI21_X1 i_4526 (.A(n_5181), .B1(inputB[5]), .B2(inputA[7]), .ZN(n_5148));
   XOR2_X1 i_4527 (.A(n_5150), .B(n_5149), .Z(n_1351));
   NAND2_X1 i_4528 (.A1(inputB[3]), .A2(inputA[9]), .ZN(n_5149));
   OAI21_X1 i_4530 (.A(n_5154), .B1(n_5234), .B2(n_5155), .ZN(n_5150));
   INV_X1 i_4531 (.A(n_5154), .ZN(n_5153));
   NAND2_X1 i_4532 (.A1(n_5234), .A2(n_5155), .ZN(n_5154));
   NAND2_X1 i_4534 (.A1(inputB[2]), .A2(inputA[10]), .ZN(n_5155));
   OAI21_X1 i_4535 (.A(n_5207), .B1(n_5217), .B2(n_5197), .ZN(n_1276));
   NAND2_X1 i_4536 (.A1(n_5227), .A2(n_5156), .ZN(n_1283));
   NAND2_X1 i_4538 (.A1(n_5222), .A2(n_5218), .ZN(n_5156));
   INV_X1 i_4539 (.A(n_5158), .ZN(n_1270));
   AOI21_X1 i_4540 (.A(n_1267), .B1(n_1266), .B2(n_5159), .ZN(n_5158));
   XNOR2_X1 i_4542 (.A(n_1261), .B(n_5161), .ZN(n_5159));
   INV_X1 i_4543 (.A(n_5161), .ZN(n_5160));
   AOI21_X1 i_4544 (.A(n_1206), .B1(n_1205), .B2(n_5283), .ZN(n_5161));
   XOR2_X1 i_4546 (.A(n_1306), .B(n_5162), .Z(n_1308));
   XOR2_X1 i_4547 (.A(n_5167), .B(n_5163), .Z(n_5162));
   NAND2_X1 i_4548 (.A1(inputB[5]), .A2(inputA[6]), .ZN(n_5163));
   NAND2_X1 i_4550 (.A1(n_5177), .A2(n_5171), .ZN(n_5167));
   INV_X1 i_4551 (.A(n_5172), .ZN(n_5171));
   AOI22_X1 i_4552 (.A1(inputB[3]), .A2(inputA[8]), .B1(inputB[4]), .B2(
      inputA[7]), .ZN(n_5172));
   NAND2_X1 i_4554 (.A1(n_5272), .A2(n_5181), .ZN(n_5177));
   AND2_X1 i_4555 (.A1(inputB[4]), .A2(inputA[8]), .ZN(n_5181));
   XNOR2_X1 i_4556 (.A(n_1311), .B(n_5187), .ZN(n_1313));
   INV_X1 i_4558 (.A(n_5187), .ZN(n_5182));
   AOI21_X1 i_4559 (.A(n_1252), .B1(n_1251), .B2(n_5251), .ZN(n_5187));
   INV_X1 i_4560 (.A(n_5192), .ZN(n_1260));
   AOI21_X1 i_4561 (.A(n_1257), .B1(n_1256), .B2(n_5240), .ZN(n_5192));
   XOR2_X1 i_4562 (.A(n_1301), .B(n_5196), .Z(n_1303));
   OAI21_X1 i_4563 (.A(n_5261), .B1(n_5264), .B2(n_5258), .ZN(n_5196));
   XOR2_X1 i_4564 (.A(n_5202), .B(n_5197), .Z(n_1275));
   NAND2_X1 i_4565 (.A1(inputB[11]), .A2(inputA[0]), .ZN(n_5197));
   NAND2_X1 i_4566 (.A1(n_5212), .A2(n_5207), .ZN(n_5202));
   NAND3_X1 i_4567 (.A1(inputB[10]), .A2(inputA[1]), .A3(n_5262), .ZN(n_5207));
   INV_X1 i_4568 (.A(n_5217), .ZN(n_5212));
   AOI21_X1 i_4569 (.A(n_5262), .B1(inputB[10]), .B2(inputA[1]), .ZN(n_5217));
   XOR2_X1 i_4570 (.A(n_5221), .B(n_5218), .Z(n_1282));
   AND2_X1 i_4571 (.A1(inputB[8]), .A2(inputA[3]), .ZN(n_5218));
   AND2_X1 i_4572 (.A1(n_5227), .A2(n_5222), .ZN(n_5221));
   NAND2_X1 i_4573 (.A1(n_5243), .A2(n_5230), .ZN(n_5222));
   NAND2_X1 i_4574 (.A1(n_5242), .A2(n_5229), .ZN(n_5227));
   INV_X1 i_4575 (.A(n_5230), .ZN(n_5229));
   NAND2_X1 i_4576 (.A1(inputB[7]), .A2(inputA[4]), .ZN(n_5230));
   XOR2_X1 i_4577 (.A(n_5233), .B(n_5232), .Z(n_1296));
   NAND2_X1 i_4578 (.A1(inputB[2]), .A2(inputA[9]), .ZN(n_5232));
   OAI21_X1 i_4579 (.A(n_5235), .B1(n_5279), .B2(n_5234), .ZN(n_5233));
   NAND2_X1 i_4580 (.A1(inputB[1]), .A2(inputA[11]), .ZN(n_5234));
   INV_X1 i_4581 (.A(n_5236), .ZN(n_5235));
   AOI22_X1 i_4582 (.A1(inputB[0]), .A2(inputA[11]), .B1(inputB[1]), .B2(
      inputA[10]), .ZN(n_5236));
   OAI22_X1 i_4583 (.A1(n_5279), .A2(n_5278), .B1(n_5276), .B2(n_5273), .ZN(
      n_1245));
   OAI22_X1 i_4584 (.A1(n_5294), .A2(n_5243), .B1(n_5245), .B2(n_5244), .ZN(
      n_1232));
   OAI21_X1 i_4585 (.A(n_5269), .B1(n_5271), .B2(n_5265), .ZN(n_1239));
   INV_X1 i_4586 (.A(n_5237), .ZN(n_1219));
   AOI21_X1 i_4587 (.A(n_1216), .B1(n_1215), .B2(n_5238), .ZN(n_5237));
   XOR2_X1 i_4588 (.A(n_1210), .B(n_5249), .Z(n_5238));
   XOR2_X1 i_4589 (.A(n_1256), .B(n_5240), .Z(n_1258));
   XNOR2_X1 i_4590 (.A(n_5245), .B(n_5241), .ZN(n_5240));
   AOI21_X1 i_4591 (.A(n_5244), .B1(n_5293), .B2(n_5242), .ZN(n_5241));
   INV_X1 i_4592 (.A(n_5243), .ZN(n_5242));
   NAND2_X1 i_4593 (.A1(inputB[6]), .A2(inputA[5]), .ZN(n_5243));
   AOI22_X1 i_4594 (.A1(inputB[5]), .A2(inputA[5]), .B1(inputB[6]), .B2(
      inputA[4]), .ZN(n_5244));
   NAND2_X1 i_4595 (.A1(inputB[7]), .A2(inputA[3]), .ZN(n_5245));
   INV_X1 i_4596 (.A(n_5248), .ZN(n_1214));
   AOI21_X1 i_4597 (.A(n_1211), .B1(n_1210), .B2(n_5249), .ZN(n_5248));
   XOR2_X1 i_4598 (.A(n_5252), .B(n_5250), .Z(n_5249));
   OAI21_X1 i_4599 (.A(n_5253), .B1(n_5257), .B2(n_5256), .ZN(n_5250));
   XOR2_X1 i_4600 (.A(n_1251), .B(n_5251), .Z(n_1253));
   OAI21_X1 i_4601 (.A(n_5253), .B1(n_5255), .B2(n_5252), .ZN(n_5251));
   NAND2_X1 i_4602 (.A1(inputB[0]), .A2(inputA[9]), .ZN(n_5252));
   NAND2_X1 i_4603 (.A1(n_5257), .A2(n_5256), .ZN(n_5253));
   NOR2_X1 i_4604 (.A1(n_5257), .A2(n_5256), .ZN(n_5255));
   AOI21_X1 i_4605 (.A(n_5354), .B1(n_5355), .B2(n_5350), .ZN(n_5256));
   AOI21_X1 i_4606 (.A(n_5363), .B1(n_5365), .B2(n_5360), .ZN(n_5257));
   XOR2_X1 i_4607 (.A(n_5259), .B(n_5258), .Z(n_1224));
   NAND2_X1 i_4608 (.A1(inputB[10]), .A2(inputA[0]), .ZN(n_5258));
   NAND2_X1 i_4609 (.A1(n_5263), .A2(n_5261), .ZN(n_5259));
   NAND2_X1 i_4610 (.A1(n_5313), .A2(n_5262), .ZN(n_5261));
   AND2_X1 i_4612 (.A1(inputB[9]), .A2(inputA[2]), .ZN(n_5262));
   INV_X1 i_4613 (.A(n_5264), .ZN(n_5263));
   AOI22_X1 i_4614 (.A1(inputB[8]), .A2(inputA[2]), .B1(inputB[9]), .B2(
      inputA[1]), .ZN(n_5264));
   XOR2_X1 i_4616 (.A(n_5266), .B(n_5265), .Z(n_1238));
   NAND2_X1 i_4617 (.A1(inputB[4]), .A2(inputA[6]), .ZN(n_5265));
   NAND2_X1 i_4618 (.A1(n_5270), .A2(n_5269), .ZN(n_5266));
   NAND3_X1 i_4620 (.A1(inputB[2]), .A2(inputA[8]), .A3(n_5272), .ZN(n_5269));
   INV_X1 i_4621 (.A(n_5271), .ZN(n_5270));
   AOI21_X1 i_4622 (.A(n_5272), .B1(inputB[2]), .B2(inputA[8]), .ZN(n_5271));
   AND2_X1 i_4624 (.A1(inputB[3]), .A2(inputA[7]), .ZN(n_5272));
   XOR2_X1 i_4625 (.A(n_5274), .B(n_5273), .Z(n_1244));
   NAND2_X1 i_4626 (.A1(inputB[1]), .A2(inputA[9]), .ZN(n_5273));
   OAI21_X1 i_4628 (.A(n_5277), .B1(n_5279), .B2(n_5278), .ZN(n_5274));
   INV_X1 i_4629 (.A(n_5277), .ZN(n_5276));
   NAND2_X1 i_4630 (.A1(n_5279), .A2(n_5278), .ZN(n_5277));
   AOI21_X1 i_4632 (.A(n_5332), .B1(n_5328), .B2(n_5318), .ZN(n_5278));
   NAND2_X1 i_4633 (.A1(inputB[0]), .A2(inputA[10]), .ZN(n_5279));
   AOI22_X1 i_4634 (.A1(n_5346), .A2(n_5317), .B1(n_5312), .B2(n_5303), .ZN(
      n_1179));
   AOI22_X1 i_4636 (.A1(n_5359), .A2(n_5294), .B1(n_5292), .B2(n_5284), .ZN(
      n_1186));
   INV_X1 i_4637 (.A(n_5282), .ZN(n_1173));
   AOI21_X1 i_4638 (.A(n_1170), .B1(n_1137), .B2(n_1169), .ZN(n_5282));
   XOR2_X1 i_4640 (.A(n_1205), .B(n_5283), .Z(n_1207));
   XOR2_X1 i_4641 (.A(n_5288), .B(n_5284), .Z(n_5283));
   NAND2_X1 i_4642 (.A1(inputB[6]), .A2(inputA[3]), .ZN(n_5284));
   OAI21_X1 i_4644 (.A(n_5292), .B1(n_5356), .B2(n_5293), .ZN(n_5288));
   NAND2_X1 i_4645 (.A1(n_5356), .A2(n_5293), .ZN(n_5292));
   INV_X1 i_4646 (.A(n_5294), .ZN(n_5293));
   NAND2_X1 i_4648 (.A1(inputB[5]), .A2(inputA[4]), .ZN(n_5294));
   INV_X1 i_4649 (.A(n_5298), .ZN(n_1168));
   AOI21_X1 i_4650 (.A(n_1165), .B1(n_1164), .B2(n_5333), .ZN(n_5298));
   INV_X1 i_4652 (.A(n_5302), .ZN(n_1163));
   AOI21_X1 i_4653 (.A(n_1160), .B1(n_1159), .B2(n_5349), .ZN(n_5302));
   XOR2_X1 i_4654 (.A(n_5308), .B(n_5303), .Z(n_1178));
   NAND2_X1 i_4656 (.A1(inputB[9]), .A2(inputA[0]), .ZN(n_5303));
   OAI21_X1 i_4657 (.A(n_5312), .B1(n_5345), .B2(n_5313), .ZN(n_5308));
   NAND2_X1 i_4658 (.A1(n_5345), .A2(n_5313), .ZN(n_5312));
   INV_X1 i_4660 (.A(n_5317), .ZN(n_5313));
   NAND2_X1 i_4661 (.A1(inputB[8]), .A2(inputA[1]), .ZN(n_5317));
   XOR2_X1 i_4662 (.A(n_5323), .B(n_5318), .Z(n_1192));
   AND2_X1 i_4664 (.A1(inputB[3]), .A2(inputA[6]), .ZN(n_5318));
   NOR2_X1 i_4665 (.A1(n_5332), .A2(n_5329), .ZN(n_5323));
   INV_X1 i_4666 (.A(n_5329), .ZN(n_5328));
   AOI21_X1 i_4667 (.A(n_5366), .B1(inputB[2]), .B2(inputA[7]), .ZN(n_5329));
   AND3_X1 i_4668 (.A1(inputB[2]), .A2(inputA[7]), .A3(n_5366), .ZN(n_5332));
   OAI21_X1 i_4669 (.A(n_5344), .B1(n_5343), .B2(n_5338), .ZN(n_1141));
   XOR2_X1 i_4670 (.A(n_1164), .B(n_5333), .Z(n_1166));
   XOR2_X1 i_4671 (.A(n_5340), .B(n_5338), .Z(n_5333));
   NAND2_X1 i_4672 (.A1(inputB[8]), .A2(inputA[0]), .ZN(n_5338));
   NAND2_X1 i_4673 (.A1(n_5344), .A2(n_5342), .ZN(n_5340));
   INV_X1 i_4674 (.A(n_5343), .ZN(n_5342));
   AOI22_X1 i_4675 (.A1(inputB[6]), .A2(inputA[2]), .B1(inputB[7]), .B2(
      inputA[1]), .ZN(n_5343));
   NAND2_X1 i_4676 (.A1(n_5386), .A2(n_5345), .ZN(n_5344));
   INV_X1 i_4677 (.A(n_5346), .ZN(n_5345));
   NAND2_X1 i_4678 (.A1(inputB[7]), .A2(inputA[2]), .ZN(n_5346));
   INV_X1 i_4679 (.A(n_5347), .ZN(n_1135));
   AOI21_X1 i_4680 (.A(n_1132), .B1(n_1103), .B2(n_1131), .ZN(n_5347));
   INV_X1 i_4681 (.A(n_5348), .ZN(n_1130));
   AOI21_X1 i_4682 (.A(n_1127), .B1(n_1126), .B2(n_5370), .ZN(n_5348));
   XOR2_X1 i_4683 (.A(n_1159), .B(n_5349), .Z(n_1161));
   OAI21_X1 i_4684 (.A(n_5376), .B1(n_5377), .B2(n_5373), .ZN(n_5349));
   XOR2_X1 i_4685 (.A(n_5352), .B(n_5350), .Z(n_1147));
   NAND2_X1 i_4686 (.A1(inputB[5]), .A2(inputA[3]), .ZN(n_5350));
   NAND2_X1 i_4687 (.A1(n_5355), .A2(n_5353), .ZN(n_5352));
   INV_X1 i_4688 (.A(n_5354), .ZN(n_5353));
   AOI22_X1 i_4689 (.A1(inputB[3]), .A2(inputA[5]), .B1(inputB[4]), .B2(
      inputA[4]), .ZN(n_5354));
   NAND2_X1 i_4690 (.A1(n_5407), .A2(n_5356), .ZN(n_5355));
   INV_X1 i_4691 (.A(n_5359), .ZN(n_5356));
   NAND2_X1 i_4692 (.A1(inputB[4]), .A2(inputA[5]), .ZN(n_5359));
   XOR2_X1 i_4693 (.A(n_5361), .B(n_5360), .Z(n_1154));
   NAND2_X1 i_4694 (.A1(inputB[2]), .A2(inputA[6]), .ZN(n_5360));
   NAND2_X1 i_4695 (.A1(n_5365), .A2(n_5362), .ZN(n_5361));
   INV_X1 i_4696 (.A(n_5363), .ZN(n_5362));
   AOI22_X1 i_4697 (.A1(inputB[0]), .A2(inputA[8]), .B1(inputB[1]), .B2(
      inputA[7]), .ZN(n_5363));
   NAND2_X1 i_4698 (.A1(n_5371), .A2(n_5366), .ZN(n_5365));
   AND2_X1 i_4699 (.A1(inputB[1]), .A2(inputA[8]), .ZN(n_5366));
   AOI22_X1 i_4700 (.A1(n_5449), .A2(n_5391), .B1(n_5385), .B2(n_5381), .ZN(
      n_1107));
   OAI21_X1 i_4701 (.A(n_5401), .B1(n_5406), .B2(n_5396), .ZN(n_1114));
   INV_X1 i_4702 (.A(n_5367), .ZN(n_1101));
   AOI21_X1 i_4703 (.A(n_1098), .B1(n_1097), .B2(n_5368), .ZN(n_5367));
   XOR2_X1 i_4704 (.A(n_5411), .B(n_5369), .Z(n_5368));
   OAI21_X1 i_4705 (.A(n_5415), .B1(n_5420), .B2(n_5417), .ZN(n_5369));
   XOR2_X1 i_4706 (.A(n_1126), .B(n_5370), .Z(n_1128));
   XOR2_X1 i_4707 (.A(n_5374), .B(n_5371), .Z(n_5370));
   INV_X1 i_4708 (.A(n_5373), .ZN(n_5371));
   NAND2_X1 i_4709 (.A1(inputB[0]), .A2(inputA[7]), .ZN(n_5373));
   NOR2_X1 i_4710 (.A1(n_5377), .A2(n_5375), .ZN(n_5374));
   INV_X1 i_4711 (.A(n_5376), .ZN(n_5375));
   NAND3_X1 i_4712 (.A1(inputB[1]), .A2(inputA[6]), .A3(n_5380), .ZN(n_5376));
   AOI21_X1 i_4713 (.A(n_5380), .B1(inputB[1]), .B2(inputA[6]), .ZN(n_5377));
   OAI21_X1 i_4714 (.A(n_5456), .B1(n_5458), .B2(n_5452), .ZN(n_5380));
   XOR2_X1 i_4715 (.A(n_5382), .B(n_5381), .Z(n_1106));
   NAND2_X1 i_4716 (.A1(inputB[7]), .A2(inputA[0]), .ZN(n_5381));
   OAI21_X1 i_4717 (.A(n_5385), .B1(n_5448), .B2(n_5386), .ZN(n_5382));
   NAND2_X1 i_4719 (.A1(n_5448), .A2(n_5386), .ZN(n_5385));
   INV_X1 i_4720 (.A(n_5391), .ZN(n_5386));
   NAND2_X1 i_4721 (.A1(inputB[6]), .A2(inputA[1]), .ZN(n_5391));
   XOR2_X1 i_4723 (.A(n_5397), .B(n_5396), .Z(n_1113));
   NAND2_X1 i_4724 (.A1(inputB[4]), .A2(inputA[3]), .ZN(n_5396));
   NAND2_X1 i_4725 (.A1(n_5405), .A2(n_5401), .ZN(n_5397));
   NAND3_X1 i_4727 (.A1(inputB[2]), .A2(inputA[5]), .A3(n_5407), .ZN(n_5401));
   INV_X1 i_4728 (.A(n_5406), .ZN(n_5405));
   AOI21_X1 i_4729 (.A(n_5407), .B1(inputB[2]), .B2(inputA[5]), .ZN(n_5406));
   AND2_X1 i_4731 (.A1(inputB[3]), .A2(inputA[4]), .ZN(n_5407));
   OAI21_X1 i_4732 (.A(n_5415), .B1(n_5416), .B2(n_5411), .ZN(n_1092));
   NAND2_X1 i_4733 (.A1(inputB[0]), .A2(inputA[6]), .ZN(n_5411));
   NAND2_X1 i_4735 (.A1(n_5420), .A2(n_5417), .ZN(n_5415));
   NOR2_X1 i_4736 (.A1(n_5420), .A2(n_5417), .ZN(n_5416));
   AOI22_X1 i_4737 (.A1(n_5472), .A2(n_5464), .B1(n_5462), .B2(n_5460), .ZN(
      n_5417));
   OAI21_X1 i_4739 (.A(n_5441), .B1(n_5436), .B2(n_5431), .ZN(n_5420));
   OAI21_X1 i_4740 (.A(n_5447), .B1(n_5451), .B2(n_5443), .ZN(n_1078));
   INV_X1 i_4741 (.A(n_5421), .ZN(n_1072));
   AOI21_X1 i_4743 (.A(n_1069), .B1(n_1068), .B2(n_5426), .ZN(n_5421));
   XOR2_X1 i_4744 (.A(n_5432), .B(n_5431), .Z(n_5426));
   NAND2_X1 i_4745 (.A1(inputB[2]), .A2(inputA[3]), .ZN(n_5431));
   NAND2_X1 i_4747 (.A1(n_5441), .A2(n_5435), .ZN(n_5432));
   INV_X1 i_4748 (.A(n_5436), .ZN(n_5435));
   AOI22_X1 i_4749 (.A1(inputB[1]), .A2(inputA[4]), .B1(inputB[0]), .B2(
      inputA[5]), .ZN(n_5436));
   NAND3_X1 i_4751 (.A1(inputB[0]), .A2(inputA[4]), .A3(n_5459), .ZN(n_5441));
   XOR2_X1 i_4752 (.A(n_5446), .B(n_5443), .Z(n_1077));
   NAND2_X1 i_4753 (.A1(inputB[6]), .A2(inputA[0]), .ZN(n_5443));
   NAND2_X1 i_4755 (.A1(n_5450), .A2(n_5447), .ZN(n_5446));
   NAND2_X1 i_4756 (.A1(n_5463), .A2(n_5448), .ZN(n_5447));
   INV_X1 i_4757 (.A(n_5449), .ZN(n_5448));
   NAND2_X1 i_4759 (.A1(inputB[5]), .A2(inputA[2]), .ZN(n_5449));
   INV_X1 i_4760 (.A(n_5451), .ZN(n_5450));
   AOI22_X1 i_4761 (.A1(inputB[4]), .A2(inputA[2]), .B1(inputB[5]), .B2(
      inputA[1]), .ZN(n_5451));
   XOR2_X1 i_4763 (.A(n_5455), .B(n_5452), .Z(n_1084));
   NAND2_X1 i_4764 (.A1(inputB[3]), .A2(inputA[3]), .ZN(n_5452));
   NAND2_X1 i_4765 (.A1(n_5457), .A2(n_5456), .ZN(n_5455));
   NAND3_X1 i_4767 (.A1(inputB[2]), .A2(inputA[4]), .A3(n_5459), .ZN(n_5456));
   INV_X1 i_4768 (.A(n_5458), .ZN(n_5457));
   AOI21_X1 i_4769 (.A(n_5459), .B1(inputB[2]), .B2(inputA[4]), .ZN(n_5458));
   AND2_X1 i_4770 (.A1(inputB[1]), .A2(inputA[5]), .ZN(n_5459));
   XOR2_X1 i_4771 (.A(n_5461), .B(n_5460), .Z(n_1056));
   NAND2_X1 i_4772 (.A1(inputB[5]), .A2(inputA[0]), .ZN(n_5460));
   OAI21_X1 i_4773 (.A(n_5462), .B1(n_5471), .B2(n_5463), .ZN(n_5461));
   NAND2_X1 i_4774 (.A1(n_5471), .A2(n_5463), .ZN(n_5462));
   INV_X1 i_4775 (.A(n_5464), .ZN(n_5463));
   NAND2_X1 i_4776 (.A1(inputB[4]), .A2(inputA[1]), .ZN(n_5464));
   AOI21_X1 i_4777 (.A(n_5469), .B1(n_5470), .B2(n_5465), .ZN(n_1040));
   NAND2_X1 i_4778 (.A1(inputB[4]), .A2(inputA[0]), .ZN(n_5465));
   INV_X1 i_4779 (.A(n_5469), .ZN(n_5466));
   AOI22_X1 i_4780 (.A1(inputB[2]), .A2(inputA[2]), .B1(inputB[3]), .B2(
      inputA[1]), .ZN(n_5469));
   NAND3_X1 i_4781 (.A1(inputB[2]), .A2(inputA[1]), .A3(n_5471), .ZN(n_5470));
   INV_X1 i_4782 (.A(n_5472), .ZN(n_5471));
   NAND2_X1 i_4783 (.A1(inputB[3]), .A2(inputA[2]), .ZN(n_5472));
   OAI22_X1 i_4784 (.A1(n_5479), .A2(n_1046), .B1(n_5495), .B2(n_5473), .ZN(
      n_1045));
   NAND2_X1 i_4785 (.A1(inputA[4]), .A2(n_5477), .ZN(n_5473));
   NOR2_X1 i_4786 (.A1(n_5478), .A2(n_5476), .ZN(n_1046));
   AOI21_X1 i_4787 (.A(n_5496), .B1(inputB[1]), .B2(inputA[4]), .ZN(n_5476));
   INV_X1 i_4788 (.A(n_5478), .ZN(n_5477));
   NAND2_X1 i_4789 (.A1(inputB[0]), .A2(inputA[3]), .ZN(n_5478));
   AOI22_X1 i_4790 (.A1(inputB[1]), .A2(inputA[3]), .B1(inputB[0]), .B2(
      inputA[4]), .ZN(n_5479));
   AOI21_X1 i_4791 (.A(n_5482), .B1(n_5483), .B2(n_5480), .ZN(n_1030));
   NAND2_X1 i_4792 (.A1(inputB[3]), .A2(inputA[0]), .ZN(n_5480));
   INV_X1 i_4793 (.A(n_5482), .ZN(n_5481));
   AOI22_X1 i_4794 (.A1(inputB[2]), .A2(inputA[1]), .B1(inputB[1]), .B2(
      inputA[2]), .ZN(n_5482));
   NAND3_X1 i_4795 (.A1(inputB[2]), .A2(inputA[2]), .A3(n_5730), .ZN(n_5483));
   AOI21_X1 i_4796 (.A(n_5484), .B1(result[0]), .B2(n_5730), .ZN(result[1]));
   AOI22_X1 i_4797 (.A1(inputB[1]), .A2(inputA[0]), .B1(inputB[0]), .B2(
      inputA[1]), .ZN(n_5484));
   XOR2_X1 i_4798 (.A(n_5490), .B(n_5485), .Z(result[2]));
   XOR2_X1 i_4799 (.A(n_5734), .B(n_5486), .Z(n_5485));
   NAND2_X1 i_4800 (.A1(result[0]), .A2(n_5730), .ZN(n_5486));
   AOI21_X1 i_4801 (.A(n_5496), .B1(n_5731), .B2(n_5729), .ZN(n_5490));
   INV_X1 i_4802 (.A(n_5496), .ZN(n_5495));
   NOR2_X1 i_4803 (.A1(n_5731), .A2(n_5729), .ZN(n_5496));
   XOR2_X1 i_4804 (.A(n_128), .B(n_5728), .Z(result[3]));
   XNOR2_X1 i_4805 (.A(n_130), .B(n_5727), .ZN(result[4]));
   XNOR2_X1 i_4806 (.A(n_132), .B(n_5725), .ZN(result[5]));
   XNOR2_X1 i_4807 (.A(n_134), .B(n_5722), .ZN(result[6]));
   XNOR2_X1 i_4808 (.A(n_136), .B(n_5715), .ZN(result[7]));
   XNOR2_X1 i_4809 (.A(n_138), .B(n_5711), .ZN(result[8]));
   XNOR2_X1 i_4810 (.A(n_140), .B(n_5706), .ZN(result[9]));
   XNOR2_X1 i_4811 (.A(n_142), .B(n_5700), .ZN(result[10]));
   XNOR2_X1 i_4812 (.A(n_144), .B(n_5696), .ZN(result[11]));
   XNOR2_X1 i_4813 (.A(n_146), .B(n_5691), .ZN(result[12]));
   XNOR2_X1 i_4814 (.A(n_148), .B(n_5685), .ZN(result[13]));
   XNOR2_X1 i_4815 (.A(n_150), .B(n_5680), .ZN(result[14]));
   XNOR2_X1 i_4816 (.A(n_152), .B(n_5675), .ZN(result[15]));
   XNOR2_X1 i_4817 (.A(n_154), .B(n_5670), .ZN(result[16]));
   XNOR2_X1 i_4818 (.A(n_156), .B(n_5667), .ZN(result[17]));
   XNOR2_X1 i_4819 (.A(n_158), .B(n_5665), .ZN(result[18]));
   XNOR2_X1 i_4820 (.A(n_160), .B(n_5663), .ZN(result[19]));
   XNOR2_X1 i_4822 (.A(n_162), .B(n_5659), .ZN(result[20]));
   XNOR2_X1 i_4823 (.A(n_164), .B(n_5657), .ZN(result[21]));
   XNOR2_X1 i_4824 (.A(n_166), .B(n_5655), .ZN(result[22]));
   XNOR2_X1 i_4826 (.A(n_168), .B(n_5652), .ZN(result[23]));
   XNOR2_X1 i_4827 (.A(n_170), .B(n_5650), .ZN(result[24]));
   XNOR2_X1 i_4828 (.A(n_172), .B(n_5648), .ZN(result[25]));
   XNOR2_X1 i_4830 (.A(n_174), .B(n_5645), .ZN(result[26]));
   XNOR2_X1 i_4831 (.A(n_176), .B(n_5643), .ZN(result[27]));
   XNOR2_X1 i_4832 (.A(n_178), .B(n_5641), .ZN(result[28]));
   XNOR2_X1 i_4834 (.A(n_180), .B(n_5639), .ZN(result[29]));
   XNOR2_X1 i_4835 (.A(n_182), .B(n_5634), .ZN(result[30]));
   XNOR2_X1 i_4836 (.A(n_184), .B(n_5628), .ZN(result[31]));
   XNOR2_X1 i_4838 (.A(n_186), .B(n_5624), .ZN(result[32]));
   XNOR2_X1 i_4839 (.A(n_188), .B(n_5615), .ZN(result[33]));
   XNOR2_X1 i_4840 (.A(n_190), .B(n_5609), .ZN(result[34]));
   XNOR2_X1 i_4842 (.A(n_192), .B(n_5604), .ZN(result[35]));
   XNOR2_X1 i_4843 (.A(n_194), .B(n_5599), .ZN(result[36]));
   XNOR2_X1 i_4844 (.A(n_196), .B(n_5594), .ZN(result[37]));
   XNOR2_X1 i_4846 (.A(n_198), .B(n_5588), .ZN(result[38]));
   XNOR2_X1 i_4847 (.A(n_200), .B(n_5584), .ZN(result[39]));
   XNOR2_X1 i_4848 (.A(n_202), .B(n_5582), .ZN(result[40]));
   XNOR2_X1 i_4850 (.A(n_204), .B(n_5578), .ZN(result[41]));
   XNOR2_X1 i_4851 (.A(n_206), .B(n_5576), .ZN(result[42]));
   XNOR2_X1 i_4852 (.A(n_208), .B(n_5573), .ZN(result[43]));
   XNOR2_X1 i_4854 (.A(n_210), .B(n_5571), .ZN(result[44]));
   XNOR2_X1 i_4855 (.A(n_212), .B(n_5569), .ZN(result[45]));
   XNOR2_X1 i_4856 (.A(n_214), .B(n_5567), .ZN(result[46]));
   XNOR2_X1 i_4858 (.A(n_216), .B(n_5564), .ZN(result[47]));
   XNOR2_X1 i_4859 (.A(n_218), .B(n_5562), .ZN(result[48]));
   XNOR2_X1 i_4860 (.A(n_220), .B(n_5558), .ZN(result[49]));
   XNOR2_X1 i_4862 (.A(n_222), .B(n_5556), .ZN(result[50]));
   XNOR2_X1 i_4863 (.A(n_224), .B(n_5554), .ZN(result[51]));
   XNOR2_X1 i_4864 (.A(n_226), .B(n_5551), .ZN(result[52]));
   XNOR2_X1 i_4866 (.A(n_228), .B(n_5549), .ZN(result[53]));
   XNOR2_X1 i_4867 (.A(n_230), .B(n_5547), .ZN(result[54]));
   XNOR2_X1 i_4868 (.A(n_232), .B(n_5545), .ZN(result[55]));
   XNOR2_X1 i_4869 (.A(n_234), .B(n_5542), .ZN(result[56]));
   XNOR2_X1 i_4870 (.A(n_236), .B(n_5535), .ZN(result[57]));
   XNOR2_X1 i_4871 (.A(n_238), .B(n_5531), .ZN(result[58]));
   XNOR2_X1 i_4872 (.A(n_240), .B(n_5525), .ZN(result[59]));
   XNOR2_X1 i_4873 (.A(n_242), .B(n_5519), .ZN(result[60]));
   XNOR2_X1 i_4874 (.A(n_244), .B(n_5511), .ZN(result[61]));
   XOR2_X1 i_4875 (.A(n_5505), .B(n_5500), .Z(result[62]));
   NAND2_X1 i_4876 (.A1(n_5737), .A2(n_5735), .ZN(n_5500));
   INV_X1 i_4877 (.A(n_5504), .ZN(result[63]));
   AOI21_X1 i_4878 (.A(n_5736), .B1(n_5737), .B2(n_5505), .ZN(n_5504));
   AOI21_X1 i_4879 (.A(n_245), .B1(n_244), .B2(n_5510), .ZN(n_5505));
   INV_X1 i_4880 (.A(n_5511), .ZN(n_5510));
   AOI21_X1 i_4881 (.A(n_243), .B1(n_242), .B2(n_5515), .ZN(n_5511));
   INV_X1 i_4882 (.A(n_5519), .ZN(n_5515));
   AOI21_X1 i_4883 (.A(n_241), .B1(n_240), .B2(n_5520), .ZN(n_5519));
   INV_X1 i_4884 (.A(n_5525), .ZN(n_5520));
   AOI21_X1 i_4885 (.A(n_239), .B1(n_238), .B2(n_5530), .ZN(n_5525));
   INV_X1 i_4886 (.A(n_5531), .ZN(n_5530));
   AOI21_X1 i_4887 (.A(n_237), .B1(n_236), .B2(n_5534), .ZN(n_5531));
   INV_X1 i_4888 (.A(n_5535), .ZN(n_5534));
   AOI21_X1 i_4889 (.A(n_235), .B1(n_234), .B2(n_5540), .ZN(n_5535));
   INV_X1 i_4890 (.A(n_5542), .ZN(n_5540));
   AOI21_X1 i_4891 (.A(n_233), .B1(n_232), .B2(n_5544), .ZN(n_5542));
   INV_X1 i_4892 (.A(n_5545), .ZN(n_5544));
   AOI21_X1 i_4893 (.A(n_231), .B1(n_230), .B2(n_5546), .ZN(n_5545));
   INV_X1 i_4894 (.A(n_5547), .ZN(n_5546));
   AOI21_X1 i_4895 (.A(n_229), .B1(n_228), .B2(n_5548), .ZN(n_5547));
   INV_X1 i_4896 (.A(n_5549), .ZN(n_5548));
   AOI21_X1 i_4897 (.A(n_227), .B1(n_226), .B2(n_5550), .ZN(n_5549));
   INV_X1 i_4898 (.A(n_5551), .ZN(n_5550));
   AOI21_X1 i_4899 (.A(n_225), .B1(n_224), .B2(n_5552), .ZN(n_5551));
   INV_X1 i_4900 (.A(n_5554), .ZN(n_5552));
   AOI21_X1 i_4901 (.A(n_223), .B1(n_222), .B2(n_5555), .ZN(n_5554));
   INV_X1 i_4902 (.A(n_5556), .ZN(n_5555));
   AOI21_X1 i_4903 (.A(n_221), .B1(n_220), .B2(n_5557), .ZN(n_5556));
   INV_X1 i_4904 (.A(n_5558), .ZN(n_5557));
   AOI21_X1 i_4905 (.A(n_219), .B1(n_218), .B2(n_5561), .ZN(n_5558));
   INV_X1 i_4906 (.A(n_5562), .ZN(n_5561));
   AOI21_X1 i_4907 (.A(n_217), .B1(n_216), .B2(n_5563), .ZN(n_5562));
   INV_X1 i_4908 (.A(n_5564), .ZN(n_5563));
   AOI21_X1 i_4909 (.A(n_215), .B1(n_214), .B2(n_5565), .ZN(n_5564));
   INV_X1 i_4910 (.A(n_5567), .ZN(n_5565));
   AOI21_X1 i_4911 (.A(n_213), .B1(n_212), .B2(n_5568), .ZN(n_5567));
   INV_X1 i_4913 (.A(n_5569), .ZN(n_5568));
   AOI21_X1 i_4914 (.A(n_211), .B1(n_210), .B2(n_5570), .ZN(n_5569));
   INV_X1 i_4915 (.A(n_5571), .ZN(n_5570));
   AOI21_X1 i_4917 (.A(n_209), .B1(n_208), .B2(n_5572), .ZN(n_5571));
   INV_X1 i_4918 (.A(n_5573), .ZN(n_5572));
   AOI21_X1 i_4919 (.A(n_207), .B1(n_206), .B2(n_5575), .ZN(n_5573));
   INV_X1 i_4921 (.A(n_5576), .ZN(n_5575));
   AOI21_X1 i_4922 (.A(n_205), .B1(n_204), .B2(n_5577), .ZN(n_5576));
   INV_X1 i_4923 (.A(n_5578), .ZN(n_5577));
   AOI21_X1 i_4925 (.A(n_203), .B1(n_202), .B2(n_5579), .ZN(n_5578));
   INV_X1 i_4926 (.A(n_5582), .ZN(n_5579));
   AOI21_X1 i_4927 (.A(n_201), .B1(n_200), .B2(n_5583), .ZN(n_5582));
   INV_X1 i_4929 (.A(n_5584), .ZN(n_5583));
   AOI21_X1 i_4930 (.A(n_199), .B1(n_198), .B2(n_5585), .ZN(n_5584));
   INV_X1 i_4931 (.A(n_5588), .ZN(n_5585));
   AOI21_X1 i_4933 (.A(n_197), .B1(n_196), .B2(n_5589), .ZN(n_5588));
   INV_X1 i_4934 (.A(n_5594), .ZN(n_5589));
   AOI21_X1 i_4935 (.A(n_195), .B1(n_194), .B2(n_5598), .ZN(n_5594));
   INV_X1 i_4937 (.A(n_5599), .ZN(n_5598));
   AOI21_X1 i_4938 (.A(n_193), .B1(n_192), .B2(n_5600), .ZN(n_5599));
   INV_X1 i_4939 (.A(n_5604), .ZN(n_5600));
   AOI21_X1 i_4941 (.A(n_191), .B1(n_190), .B2(n_5608), .ZN(n_5604));
   INV_X1 i_4942 (.A(n_5609), .ZN(n_5608));
   AOI21_X1 i_4943 (.A(n_189), .B1(n_188), .B2(n_5614), .ZN(n_5609));
   INV_X1 i_4945 (.A(n_5615), .ZN(n_5614));
   AOI21_X1 i_4946 (.A(n_187), .B1(n_186), .B2(n_5619), .ZN(n_5615));
   INV_X1 i_4947 (.A(n_5624), .ZN(n_5619));
   AOI21_X1 i_4949 (.A(n_185), .B1(n_184), .B2(n_5625), .ZN(n_5624));
   INV_X1 i_4950 (.A(n_5628), .ZN(n_5625));
   AOI21_X1 i_4951 (.A(n_183), .B1(n_182), .B2(n_5629), .ZN(n_5628));
   INV_X1 i_4953 (.A(n_5634), .ZN(n_5629));
   AOI21_X1 i_4954 (.A(n_181), .B1(n_180), .B2(n_5636), .ZN(n_5634));
   INV_X1 i_4955 (.A(n_5639), .ZN(n_5636));
   AOI21_X1 i_4957 (.A(n_179), .B1(n_178), .B2(n_5640), .ZN(n_5639));
   INV_X1 i_4958 (.A(n_5641), .ZN(n_5640));
   AOI21_X1 i_4959 (.A(n_177), .B1(n_176), .B2(n_5642), .ZN(n_5641));
   INV_X1 i_4960 (.A(n_5643), .ZN(n_5642));
   AOI21_X1 i_4961 (.A(n_175), .B1(n_174), .B2(n_5644), .ZN(n_5643));
   INV_X1 i_4962 (.A(n_5645), .ZN(n_5644));
   AOI21_X1 i_4963 (.A(n_173), .B1(n_172), .B2(n_5646), .ZN(n_5645));
   INV_X1 i_4964 (.A(n_5648), .ZN(n_5646));
   AOI21_X1 i_4965 (.A(n_171), .B1(n_170), .B2(n_5649), .ZN(n_5648));
   INV_X1 i_4966 (.A(n_5650), .ZN(n_5649));
   AOI21_X1 i_4967 (.A(n_169), .B1(n_168), .B2(n_5651), .ZN(n_5650));
   INV_X1 i_4968 (.A(n_5652), .ZN(n_5651));
   AOI21_X1 i_4969 (.A(n_167), .B1(n_166), .B2(n_5654), .ZN(n_5652));
   INV_X1 i_4970 (.A(n_5655), .ZN(n_5654));
   AOI21_X1 i_4971 (.A(n_165), .B1(n_164), .B2(n_5656), .ZN(n_5655));
   INV_X1 i_4972 (.A(n_5657), .ZN(n_5656));
   AOI21_X1 i_4973 (.A(n_163), .B1(n_162), .B2(n_5658), .ZN(n_5657));
   INV_X1 i_4974 (.A(n_5659), .ZN(n_5658));
   AOI21_X1 i_4975 (.A(n_161), .B1(n_160), .B2(n_5662), .ZN(n_5659));
   INV_X1 i_4976 (.A(n_5663), .ZN(n_5662));
   AOI21_X1 i_4977 (.A(n_159), .B1(n_158), .B2(n_5664), .ZN(n_5663));
   INV_X1 i_4978 (.A(n_5665), .ZN(n_5664));
   AOI21_X1 i_4979 (.A(n_157), .B1(n_156), .B2(n_5666), .ZN(n_5665));
   INV_X1 i_4980 (.A(n_5667), .ZN(n_5666));
   AOI21_X1 i_4981 (.A(n_155), .B1(n_154), .B2(n_5669), .ZN(n_5667));
   INV_X1 i_4982 (.A(n_5670), .ZN(n_5669));
   AOI21_X1 i_4983 (.A(n_153), .B1(n_152), .B2(n_5671), .ZN(n_5670));
   INV_X1 i_4984 (.A(n_5675), .ZN(n_5671));
   AOI21_X1 i_4985 (.A(n_151), .B1(n_150), .B2(n_5679), .ZN(n_5675));
   INV_X1 i_4986 (.A(n_5680), .ZN(n_5679));
   AOI21_X1 i_4987 (.A(n_149), .B1(n_148), .B2(n_5681), .ZN(n_5680));
   INV_X1 i_4988 (.A(n_5685), .ZN(n_5681));
   AOI21_X1 i_4989 (.A(n_147), .B1(n_146), .B2(n_5690), .ZN(n_5685));
   INV_X1 i_4990 (.A(n_5691), .ZN(n_5690));
   AOI21_X1 i_4991 (.A(n_145), .B1(n_144), .B2(n_5695), .ZN(n_5691));
   INV_X1 i_4992 (.A(n_5696), .ZN(n_5695));
   AOI21_X1 i_4993 (.A(n_143), .B1(n_142), .B2(n_5699), .ZN(n_5696));
   INV_X1 i_4994 (.A(n_5700), .ZN(n_5699));
   AOI21_X1 i_4995 (.A(n_141), .B1(n_140), .B2(n_5705), .ZN(n_5700));
   INV_X1 i_4996 (.A(n_5706), .ZN(n_5705));
   AOI21_X1 i_4997 (.A(n_139), .B1(n_138), .B2(n_5710), .ZN(n_5706));
   INV_X1 i_4998 (.A(n_5711), .ZN(n_5710));
   AOI21_X1 i_4999 (.A(n_137), .B1(n_136), .B2(n_5714), .ZN(n_5711));
   INV_X1 i_5000 (.A(n_5715), .ZN(n_5714));
   AOI21_X1 i_5001 (.A(n_135), .B1(n_134), .B2(n_5720), .ZN(n_5715));
   INV_X1 i_5002 (.A(n_5722), .ZN(n_5720));
   AOI21_X1 i_5003 (.A(n_133), .B1(n_132), .B2(n_5723), .ZN(n_5722));
   INV_X1 i_5005 (.A(n_5725), .ZN(n_5723));
   AOI21_X1 i_5006 (.A(n_131), .B1(n_130), .B2(n_5726), .ZN(n_5725));
   INV_X1 i_5007 (.A(n_5727), .ZN(n_5726));
   AOI21_X1 i_5009 (.A(n_129), .B1(n_128), .B2(n_5728), .ZN(n_5727));
   AOI22_X1 i_5010 (.A1(n_5734), .A2(n_5733), .B1(n_5731), .B2(n_5729), .ZN(
      n_5728));
   NAND2_X1 i_5011 (.A1(inputB[2]), .A2(inputA[0]), .ZN(n_5729));
   INV_X1 i_5013 (.A(n_5731), .ZN(n_5730));
   NAND2_X1 i_5014 (.A1(inputB[1]), .A2(inputA[1]), .ZN(n_5731));
   NAND2_X1 i_5015 (.A1(n_5755), .A2(result[0]), .ZN(n_5733));
   AND2_X1 i_5017 (.A1(inputB[0]), .A2(inputA[0]), .ZN(result[0]));
   NAND2_X1 i_5018 (.A1(inputB[0]), .A2(inputA[2]), .ZN(n_5734));
   INV_X1 i_5019 (.A(n_5736), .ZN(n_5735));
   AOI21_X1 i_5021 (.A(n_5738), .B1(inputB[31]), .B2(inputA[31]), .ZN(n_5736));
   NAND3_X1 i_5022 (.A1(inputB[31]), .A2(inputA[31]), .A3(n_5738), .ZN(n_5737));
   INV_X1 i_5023 (.A(n_5741), .ZN(n_5738));
   AOI21_X1 i_5025 (.A(n_127), .B1(n_126), .B2(n_5742), .ZN(n_5741));
   AOI21_X1 i_5026 (.A(n_5746), .B1(n_5744), .B2(n_5743), .ZN(n_5742));
   AOI21_X1 i_5027 (.A(n_5746), .B1(n_5749), .B2(n_5748), .ZN(n_5743));
   INV_X1 i_5029 (.A(n_5745), .ZN(n_5744));
   NAND2_X1 i_5030 (.A1(inputB[31]), .A2(inputA[29]), .ZN(n_5745));
   NOR2_X1 i_5031 (.A1(n_5749), .A2(n_5748), .ZN(n_5746));
   AND2_X1 i_5033 (.A1(inputB[30]), .A2(inputA[30]), .ZN(n_5748));
   NAND2_X1 i_5034 (.A1(inputB[29]), .A2(inputA[31]), .ZN(n_5749));
   INV_X1 i_5035 (.A(inputA[29]), .ZN(n_5750));
   INV_X1 i_5037 (.A(inputA[30]), .ZN(n_5751));
   INV_X1 i_5038 (.A(inputA[31]), .ZN(n_5753));
   INV_X1 i_5039 (.A(inputB[1]), .ZN(n_5754));
   INV_X1 i_5041 (.A(inputB[2]), .ZN(n_5755));
   INV_X1 i_5042 (.A(inputB[3]), .ZN(n_5756));
   INV_X1 i_5043 (.A(inputB[9]), .ZN(n_5757));
   INV_X1 i_5045 (.A(inputB[11]), .ZN(n_5758));
   INV_X1 i_5046 (.A(inputB[17]), .ZN(n_5762));
   INV_X1 i_5047 (.A(inputB[24]), .ZN(n_5767));
endmodule

module multiplyTimes(inputA, inputB, result);
   input [31:0]inputA;
   input [31:0]inputB;
   output [63:0]result;

   datapath i_0 (.inputB(inputB), .inputA(inputA), .result(result));
endmodule

module registerNbits__2_2(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits__2_5(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits__2_8(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module integrationMult(clk, reset, en, inputA, inputB, result);
   input clk;
   input reset;
   input en;
   input [31:0]inputA;
   input [31:0]inputB;
   output [63:0]result;

   wire [31:0]outB_reg;
   wire [31:0]outA_reg;
   wire [31:0]A_reg;
   wire [31:0]B_reg;

   multiplyTimes mult (.inputA(A_reg), .inputB(B_reg), .result({outA_reg[31], 
      outA_reg[30], outA_reg[29], outA_reg[28], outA_reg[27], outA_reg[26], 
      outA_reg[25], outA_reg[24], outA_reg[23], outA_reg[22], outA_reg[21], 
      outA_reg[20], outA_reg[19], outA_reg[18], outA_reg[17], outA_reg[16], 
      outA_reg[15], outA_reg[14], outA_reg[13], outA_reg[12], outA_reg[11], 
      outA_reg[10], outA_reg[9], outA_reg[8], outA_reg[7], outA_reg[6], 
      outA_reg[5], outA_reg[4], outA_reg[3], outA_reg[2], outA_reg[1], 
      outA_reg[0], outB_reg[31], outB_reg[30], outB_reg[29], outB_reg[28], 
      outB_reg[27], outB_reg[26], outB_reg[25], outB_reg[24], outB_reg[23], 
      outB_reg[22], outB_reg[21], outB_reg[20], outB_reg[19], outB_reg[18], 
      outB_reg[17], outB_reg[16], outB_reg[15], outB_reg[14], outB_reg[13], 
      outB_reg[12], outB_reg[11], outB_reg[10], outB_reg[9], outB_reg[8], 
      outB_reg[7], outB_reg[6], outB_reg[5], outB_reg[4], outB_reg[3], 
      outB_reg[2], outB_reg[1], outB_reg[0]}));
   registerNbits__2_2 regA (.clk(clk), .reset(reset), .en(en), .inp(inputA), 
      .out(A_reg));
   registerNbits__2_5 regB (.clk(clk), .reset(reset), .en(en), .inp(inputB), 
      .out(B_reg));
   registerNbits__2_8 outB (.clk(clk), .reset(reset), .en(en), .inp(outA_reg), 
      .out({result[63], result[62], result[61], result[60], result[59], 
      result[58], result[57], result[56], result[55], result[54], result[53], 
      result[52], result[51], result[50], result[49], result[48], result[47], 
      result[46], result[45], result[44], result[43], result[42], result[41], 
      result[40], result[39], result[38], result[37], result[36], result[35], 
      result[34], result[33], result[32]}));
   registerNbits outA (.clk(clk), .reset(reset), .en(en), .inp(outB_reg), 
      .out({result[31], result[30], result[29], result[28], result[27], 
      result[26], result[25], result[24], result[23], result[22], result[21], 
      result[20], result[19], result[18], result[17], result[16], result[15], 
      result[14], result[13], result[12], result[11], result[10], result[9], 
      result[8], result[7], result[6], result[5], result[4], result[3], 
      result[2], result[1], result[0]}));
endmodule
