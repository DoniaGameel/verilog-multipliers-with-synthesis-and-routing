/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Jan  3 22:44:10 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3705530235 */

module registerNbits__0_16(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits__parameterized0(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [63:0]inp;
   output [63:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[63]  (.D(n_65), .CK(n_0), .Q(out[63]), .QN());
   DFF_X1 \out_reg[62]  (.D(n_64), .CK(n_0), .Q(out[62]), .QN());
   DFF_X1 \out_reg[61]  (.D(n_63), .CK(n_0), .Q(out[61]), .QN());
   DFF_X1 \out_reg[60]  (.D(n_62), .CK(n_0), .Q(out[60]), .QN());
   DFF_X1 \out_reg[59]  (.D(n_61), .CK(n_0), .Q(out[59]), .QN());
   DFF_X1 \out_reg[58]  (.D(n_60), .CK(n_0), .Q(out[58]), .QN());
   DFF_X1 \out_reg[57]  (.D(n_59), .CK(n_0), .Q(out[57]), .QN());
   DFF_X1 \out_reg[56]  (.D(n_58), .CK(n_0), .Q(out[56]), .QN());
   DFF_X1 \out_reg[55]  (.D(n_57), .CK(n_0), .Q(out[55]), .QN());
   DFF_X1 \out_reg[54]  (.D(n_56), .CK(n_0), .Q(out[54]), .QN());
   DFF_X1 \out_reg[53]  (.D(n_55), .CK(n_0), .Q(out[53]), .QN());
   DFF_X1 \out_reg[52]  (.D(n_54), .CK(n_0), .Q(out[52]), .QN());
   DFF_X1 \out_reg[51]  (.D(n_53), .CK(n_0), .Q(out[51]), .QN());
   DFF_X1 \out_reg[50]  (.D(n_52), .CK(n_0), .Q(out[50]), .QN());
   DFF_X1 \out_reg[49]  (.D(n_51), .CK(n_0), .Q(out[49]), .QN());
   DFF_X1 \out_reg[48]  (.D(n_50), .CK(n_0), .Q(out[48]), .QN());
   DFF_X1 \out_reg[47]  (.D(n_49), .CK(n_0), .Q(out[47]), .QN());
   DFF_X1 \out_reg[46]  (.D(n_48), .CK(n_0), .Q(out[46]), .QN());
   DFF_X1 \out_reg[45]  (.D(n_47), .CK(n_0), .Q(out[45]), .QN());
   DFF_X1 \out_reg[44]  (.D(n_46), .CK(n_0), .Q(out[44]), .QN());
   DFF_X1 \out_reg[43]  (.D(n_45), .CK(n_0), .Q(out[43]), .QN());
   DFF_X1 \out_reg[42]  (.D(n_44), .CK(n_0), .Q(out[42]), .QN());
   DFF_X1 \out_reg[41]  (.D(n_43), .CK(n_0), .Q(out[41]), .QN());
   DFF_X1 \out_reg[40]  (.D(n_42), .CK(n_0), .Q(out[40]), .QN());
   DFF_X1 \out_reg[39]  (.D(n_41), .CK(n_0), .Q(out[39]), .QN());
   DFF_X1 \out_reg[38]  (.D(n_40), .CK(n_0), .Q(out[38]), .QN());
   DFF_X1 \out_reg[37]  (.D(n_39), .CK(n_0), .Q(out[37]), .QN());
   DFF_X1 \out_reg[36]  (.D(n_38), .CK(n_0), .Q(out[36]), .QN());
   DFF_X1 \out_reg[35]  (.D(n_37), .CK(n_0), .Q(out[35]), .QN());
   DFF_X1 \out_reg[34]  (.D(n_36), .CK(n_0), .Q(out[34]), .QN());
   DFF_X1 \out_reg[33]  (.D(n_35), .CK(n_0), .Q(out[33]), .QN());
   DFF_X1 \out_reg[32]  (.D(n_34), .CK(n_0), .Q(out[32]), .QN());
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
   AND2_X1 i_0_34 (.A1(n_0_0), .A2(inp[32]), .ZN(n_34));
   AND2_X1 i_0_35 (.A1(n_0_0), .A2(inp[33]), .ZN(n_35));
   AND2_X1 i_0_36 (.A1(n_0_0), .A2(inp[34]), .ZN(n_36));
   AND2_X1 i_0_37 (.A1(n_0_0), .A2(inp[35]), .ZN(n_37));
   AND2_X1 i_0_38 (.A1(n_0_0), .A2(inp[36]), .ZN(n_38));
   AND2_X1 i_0_39 (.A1(n_0_0), .A2(inp[37]), .ZN(n_39));
   AND2_X1 i_0_40 (.A1(n_0_0), .A2(inp[38]), .ZN(n_40));
   AND2_X1 i_0_41 (.A1(n_0_0), .A2(inp[39]), .ZN(n_41));
   AND2_X1 i_0_42 (.A1(n_0_0), .A2(inp[40]), .ZN(n_42));
   AND2_X1 i_0_43 (.A1(n_0_0), .A2(inp[41]), .ZN(n_43));
   AND2_X1 i_0_44 (.A1(n_0_0), .A2(inp[42]), .ZN(n_44));
   AND2_X1 i_0_45 (.A1(n_0_0), .A2(inp[43]), .ZN(n_45));
   AND2_X1 i_0_46 (.A1(n_0_0), .A2(inp[44]), .ZN(n_46));
   AND2_X1 i_0_47 (.A1(n_0_0), .A2(inp[45]), .ZN(n_47));
   AND2_X1 i_0_48 (.A1(n_0_0), .A2(inp[46]), .ZN(n_48));
   AND2_X1 i_0_49 (.A1(n_0_0), .A2(inp[47]), .ZN(n_49));
   AND2_X1 i_0_50 (.A1(n_0_0), .A2(inp[48]), .ZN(n_50));
   AND2_X1 i_0_51 (.A1(n_0_0), .A2(inp[49]), .ZN(n_51));
   AND2_X1 i_0_52 (.A1(n_0_0), .A2(inp[50]), .ZN(n_52));
   AND2_X1 i_0_53 (.A1(n_0_0), .A2(inp[51]), .ZN(n_53));
   AND2_X1 i_0_54 (.A1(n_0_0), .A2(inp[52]), .ZN(n_54));
   AND2_X1 i_0_55 (.A1(n_0_0), .A2(inp[53]), .ZN(n_55));
   AND2_X1 i_0_56 (.A1(n_0_0), .A2(inp[54]), .ZN(n_56));
   AND2_X1 i_0_57 (.A1(n_0_0), .A2(inp[55]), .ZN(n_57));
   AND2_X1 i_0_58 (.A1(n_0_0), .A2(inp[56]), .ZN(n_58));
   AND2_X1 i_0_59 (.A1(n_0_0), .A2(inp[57]), .ZN(n_59));
   AND2_X1 i_0_60 (.A1(n_0_0), .A2(inp[58]), .ZN(n_60));
   AND2_X1 i_0_61 (.A1(n_0_0), .A2(inp[59]), .ZN(n_61));
   AND2_X1 i_0_62 (.A1(n_0_0), .A2(inp[60]), .ZN(n_62));
   AND2_X1 i_0_63 (.A1(n_0_0), .A2(inp[61]), .ZN(n_63));
   AND2_X1 i_0_64 (.A1(n_0_0), .A2(inp[62]), .ZN(n_64));
   AND2_X1 i_0_65 (.A1(n_0_0), .A2(inp[63]), .ZN(n_65));
endmodule

module datapath(p_0, A_reg);
   output [31:0]p_0;
   input [31:0]A_reg;

   XOR2_X1 i_0 (.A(A_reg[1]), .B(A_reg[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(A_reg[2]), .B1(A_reg[1]), .B2(A_reg[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(A_reg[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(A_reg[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(A_reg[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(A_reg[6]), .B1(n_27), .B2(A_reg[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(A_reg[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(A_reg[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(A_reg[9]), .B1(n_25), .B2(A_reg[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(A_reg[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(A_reg[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(A_reg[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(A_reg[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(A_reg[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(A_reg[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(A_reg[16]), .B1(n_19), .B2(A_reg[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(A_reg[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(A_reg[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(A_reg[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(A_reg[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(A_reg[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(A_reg[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(A_reg[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(A_reg[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(A_reg[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(A_reg[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(A_reg[27]), .B1(n_9), .B2(A_reg[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(A_reg[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(A_reg[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(A_reg[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(A_reg[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(A_reg[28]), .A3(A_reg[29]), .A4(A_reg[30]), 
      .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(A_reg[28]), .A3(A_reg[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(A_reg[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(A_reg[26]), .A3(A_reg[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(A_reg[23]), .A3(A_reg[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(A_reg[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(A_reg[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(A_reg[18]), .A3(A_reg[19]), .A4(A_reg[20]), 
      .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(A_reg[18]), .A3(A_reg[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(A_reg[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(A_reg[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(A_reg[15]), .A3(A_reg[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(A_reg[12]), .A3(A_reg[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(A_reg[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(A_reg[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(A_reg[8]), .A3(A_reg[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(A_reg[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(A_reg[5]), .A3(A_reg[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(A_reg[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(A_reg[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(A_reg[2]), .A2(A_reg[1]), .A3(A_reg[0]), .ZN(n_29));
   INV_X1 i_61 (.A(A_reg[11]), .ZN(n_30));
   INV_X1 i_62 (.A(A_reg[14]), .ZN(n_31));
   INV_X1 i_63 (.A(A_reg[21]), .ZN(n_32));
   INV_X1 i_64 (.A(A_reg[25]), .ZN(n_33));
endmodule

module datapath__0_12(partialProd, Acc, p_0);
   input [63:0]partialProd;
   input [63:0]Acc;
   output [63:0]p_0;

   HA_X1 i_0 (.A(partialProd[0]), .B(Acc[0]), .CO(n_0), .S(p_0[0]));
   HA_X1 i_1 (.A(partialProd[1]), .B(Acc[1]), .CO(n_2), .S(n_1));
   HA_X1 i_5 (.A(partialProd[2]), .B(Acc[2]), .CO(n_6), .S(n_5));
   HA_X1 i_9 (.A(partialProd[3]), .B(Acc[3]), .CO(n_10), .S(n_9));
   HA_X1 i_13 (.A(partialProd[4]), .B(Acc[4]), .CO(n_14), .S(n_13));
   HA_X1 i_17 (.A(partialProd[5]), .B(Acc[5]), .CO(n_18), .S(n_17));
   HA_X1 i_21 (.A(partialProd[6]), .B(Acc[6]), .CO(n_22), .S(n_21));
   HA_X1 i_25 (.A(partialProd[7]), .B(Acc[7]), .CO(n_26), .S(n_25));
   HA_X1 i_29 (.A(partialProd[8]), .B(Acc[8]), .CO(n_30), .S(n_29));
   HA_X1 i_33 (.A(partialProd[9]), .B(Acc[9]), .CO(n_34), .S(n_33));
   HA_X1 i_37 (.A(partialProd[10]), .B(Acc[10]), .CO(n_38), .S(n_37));
   HA_X1 i_41 (.A(partialProd[11]), .B(Acc[11]), .CO(n_42), .S(n_41));
   HA_X1 i_45 (.A(partialProd[12]), .B(Acc[12]), .CO(n_46), .S(n_45));
   HA_X1 i_49 (.A(partialProd[13]), .B(Acc[13]), .CO(n_50), .S(n_49));
   HA_X1 i_53 (.A(partialProd[14]), .B(Acc[14]), .CO(n_54), .S(n_53));
   HA_X1 i_57 (.A(partialProd[15]), .B(Acc[15]), .CO(n_58), .S(n_57));
   HA_X1 i_61 (.A(partialProd[16]), .B(Acc[16]), .CO(n_62), .S(n_61));
   HA_X1 i_65 (.A(partialProd[17]), .B(Acc[17]), .CO(n_66), .S(n_65));
   HA_X1 i_69 (.A(partialProd[18]), .B(Acc[18]), .CO(n_70), .S(n_69));
   HA_X1 i_73 (.A(partialProd[19]), .B(Acc[19]), .CO(n_74), .S(n_73));
   HA_X1 i_77 (.A(partialProd[20]), .B(Acc[20]), .CO(n_78), .S(n_77));
   HA_X1 i_81 (.A(partialProd[21]), .B(Acc[21]), .CO(n_82), .S(n_81));
   HA_X1 i_85 (.A(partialProd[22]), .B(Acc[22]), .CO(n_86), .S(n_85));
   HA_X1 i_89 (.A(partialProd[23]), .B(Acc[23]), .CO(n_90), .S(n_89));
   HA_X1 i_93 (.A(partialProd[24]), .B(Acc[24]), .CO(n_94), .S(n_93));
   HA_X1 i_97 (.A(partialProd[25]), .B(Acc[25]), .CO(n_98), .S(n_97));
   HA_X1 i_101 (.A(partialProd[26]), .B(Acc[26]), .CO(n_102), .S(n_101));
   HA_X1 i_105 (.A(partialProd[27]), .B(Acc[27]), .CO(n_106), .S(n_105));
   HA_X1 i_109 (.A(partialProd[28]), .B(Acc[28]), .CO(n_110), .S(n_109));
   HA_X1 i_113 (.A(partialProd[29]), .B(Acc[29]), .CO(n_114), .S(n_113));
   HA_X1 i_117 (.A(partialProd[30]), .B(Acc[30]), .CO(n_118), .S(n_117));
   HA_X1 i_121 (.A(partialProd[31]), .B(Acc[31]), .CO(n_122), .S(n_121));
   HA_X1 i_125 (.A(partialProd[32]), .B(Acc[32]), .CO(n_126), .S(n_125));
   HA_X1 i_129 (.A(partialProd[33]), .B(Acc[33]), .CO(n_130), .S(n_129));
   HA_X1 i_133 (.A(partialProd[34]), .B(Acc[34]), .CO(n_134), .S(n_133));
   HA_X1 i_137 (.A(partialProd[35]), .B(Acc[35]), .CO(n_138), .S(n_137));
   HA_X1 i_141 (.A(partialProd[36]), .B(Acc[36]), .CO(n_142), .S(n_141));
   HA_X1 i_145 (.A(partialProd[37]), .B(Acc[37]), .CO(n_146), .S(n_145));
   HA_X1 i_149 (.A(partialProd[38]), .B(Acc[38]), .CO(n_150), .S(n_149));
   HA_X1 i_153 (.A(partialProd[39]), .B(Acc[39]), .CO(n_154), .S(n_153));
   HA_X1 i_157 (.A(partialProd[40]), .B(Acc[40]), .CO(n_158), .S(n_157));
   HA_X1 i_161 (.A(partialProd[41]), .B(Acc[41]), .CO(n_162), .S(n_161));
   HA_X1 i_165 (.A(partialProd[42]), .B(Acc[42]), .CO(n_166), .S(n_165));
   HA_X1 i_169 (.A(partialProd[43]), .B(Acc[43]), .CO(n_170), .S(n_169));
   HA_X1 i_173 (.A(partialProd[44]), .B(Acc[44]), .CO(n_174), .S(n_173));
   HA_X1 i_177 (.A(partialProd[45]), .B(Acc[45]), .CO(n_178), .S(n_177));
   HA_X1 i_181 (.A(partialProd[46]), .B(Acc[46]), .CO(n_182), .S(n_181));
   HA_X1 i_185 (.A(partialProd[47]), .B(Acc[47]), .CO(n_186), .S(n_185));
   HA_X1 i_189 (.A(partialProd[48]), .B(Acc[48]), .CO(n_190), .S(n_189));
   HA_X1 i_193 (.A(partialProd[49]), .B(Acc[49]), .CO(n_194), .S(n_193));
   HA_X1 i_197 (.A(partialProd[50]), .B(Acc[50]), .CO(n_198), .S(n_197));
   HA_X1 i_201 (.A(partialProd[51]), .B(Acc[51]), .CO(n_202), .S(n_201));
   HA_X1 i_205 (.A(partialProd[52]), .B(Acc[52]), .CO(n_206), .S(n_205));
   HA_X1 i_209 (.A(partialProd[53]), .B(Acc[53]), .CO(n_210), .S(n_209));
   HA_X1 i_213 (.A(partialProd[54]), .B(Acc[54]), .CO(n_214), .S(n_213));
   HA_X1 i_217 (.A(partialProd[55]), .B(Acc[55]), .CO(n_218), .S(n_217));
   HA_X1 i_221 (.A(partialProd[56]), .B(Acc[56]), .CO(n_222), .S(n_221));
   HA_X1 i_225 (.A(partialProd[57]), .B(Acc[57]), .CO(n_226), .S(n_225));
   HA_X1 i_229 (.A(partialProd[58]), .B(Acc[58]), .CO(n_230), .S(n_229));
   HA_X1 i_233 (.A(partialProd[59]), .B(Acc[59]), .CO(n_234), .S(n_233));
   HA_X1 i_237 (.A(partialProd[60]), .B(Acc[60]), .CO(n_238), .S(n_237));
   HA_X1 i_241 (.A(partialProd[61]), .B(Acc[61]), .CO(n_242), .S(n_241));
   HA_X1 i_245 (.A(partialProd[62]), .B(Acc[62]), .CO(n_246), .S(n_245));
   XOR2_X1 i_2 (.A(n_0), .B(n_1), .Z(p_0[1]));
   XNOR2_X1 i_3 (.A(n_5), .B(n_248), .ZN(p_0[2]));
   XNOR2_X1 i_4 (.A(n_9), .B(n_244), .ZN(p_0[3]));
   XNOR2_X1 i_6 (.A(n_13), .B(n_240), .ZN(p_0[4]));
   XNOR2_X1 i_7 (.A(n_17), .B(n_236), .ZN(p_0[5]));
   XNOR2_X1 i_8 (.A(n_21), .B(n_232), .ZN(p_0[6]));
   XNOR2_X1 i_10 (.A(n_25), .B(n_228), .ZN(p_0[7]));
   XNOR2_X1 i_11 (.A(n_29), .B(n_224), .ZN(p_0[8]));
   XNOR2_X1 i_12 (.A(n_33), .B(n_220), .ZN(p_0[9]));
   XNOR2_X1 i_14 (.A(n_37), .B(n_216), .ZN(p_0[10]));
   XNOR2_X1 i_15 (.A(n_41), .B(n_212), .ZN(p_0[11]));
   XNOR2_X1 i_16 (.A(n_45), .B(n_208), .ZN(p_0[12]));
   XNOR2_X1 i_18 (.A(n_49), .B(n_204), .ZN(p_0[13]));
   XNOR2_X1 i_19 (.A(n_53), .B(n_200), .ZN(p_0[14]));
   XNOR2_X1 i_20 (.A(n_57), .B(n_196), .ZN(p_0[15]));
   XNOR2_X1 i_22 (.A(n_61), .B(n_192), .ZN(p_0[16]));
   XNOR2_X1 i_23 (.A(n_65), .B(n_188), .ZN(p_0[17]));
   XNOR2_X1 i_24 (.A(n_69), .B(n_184), .ZN(p_0[18]));
   XNOR2_X1 i_26 (.A(n_73), .B(n_180), .ZN(p_0[19]));
   XNOR2_X1 i_27 (.A(n_77), .B(n_176), .ZN(p_0[20]));
   XNOR2_X1 i_28 (.A(n_81), .B(n_172), .ZN(p_0[21]));
   XNOR2_X1 i_30 (.A(n_85), .B(n_168), .ZN(p_0[22]));
   XNOR2_X1 i_31 (.A(n_89), .B(n_164), .ZN(p_0[23]));
   XNOR2_X1 i_32 (.A(n_93), .B(n_160), .ZN(p_0[24]));
   XNOR2_X1 i_34 (.A(n_97), .B(n_156), .ZN(p_0[25]));
   XNOR2_X1 i_35 (.A(n_101), .B(n_152), .ZN(p_0[26]));
   XNOR2_X1 i_36 (.A(n_105), .B(n_148), .ZN(p_0[27]));
   XNOR2_X1 i_38 (.A(n_109), .B(n_144), .ZN(p_0[28]));
   XNOR2_X1 i_39 (.A(n_113), .B(n_140), .ZN(p_0[29]));
   XNOR2_X1 i_40 (.A(n_117), .B(n_136), .ZN(p_0[30]));
   XNOR2_X1 i_42 (.A(n_121), .B(n_132), .ZN(p_0[31]));
   XNOR2_X1 i_43 (.A(n_125), .B(n_128), .ZN(p_0[32]));
   XNOR2_X1 i_44 (.A(n_129), .B(n_124), .ZN(p_0[33]));
   XNOR2_X1 i_46 (.A(n_133), .B(n_120), .ZN(p_0[34]));
   XNOR2_X1 i_47 (.A(n_137), .B(n_116), .ZN(p_0[35]));
   XNOR2_X1 i_48 (.A(n_141), .B(n_112), .ZN(p_0[36]));
   XNOR2_X1 i_50 (.A(n_145), .B(n_108), .ZN(p_0[37]));
   XNOR2_X1 i_51 (.A(n_149), .B(n_104), .ZN(p_0[38]));
   XNOR2_X1 i_52 (.A(n_153), .B(n_100), .ZN(p_0[39]));
   XNOR2_X1 i_54 (.A(n_157), .B(n_96), .ZN(p_0[40]));
   XNOR2_X1 i_55 (.A(n_161), .B(n_92), .ZN(p_0[41]));
   XNOR2_X1 i_56 (.A(n_165), .B(n_88), .ZN(p_0[42]));
   XNOR2_X1 i_58 (.A(n_169), .B(n_84), .ZN(p_0[43]));
   XNOR2_X1 i_59 (.A(n_173), .B(n_80), .ZN(p_0[44]));
   XNOR2_X1 i_60 (.A(n_177), .B(n_76), .ZN(p_0[45]));
   XNOR2_X1 i_62 (.A(n_181), .B(n_72), .ZN(p_0[46]));
   XNOR2_X1 i_63 (.A(n_185), .B(n_68), .ZN(p_0[47]));
   XNOR2_X1 i_64 (.A(n_189), .B(n_64), .ZN(p_0[48]));
   XNOR2_X1 i_66 (.A(n_193), .B(n_60), .ZN(p_0[49]));
   XNOR2_X1 i_67 (.A(n_197), .B(n_56), .ZN(p_0[50]));
   XNOR2_X1 i_68 (.A(n_201), .B(n_52), .ZN(p_0[51]));
   XNOR2_X1 i_70 (.A(n_205), .B(n_48), .ZN(p_0[52]));
   XNOR2_X1 i_71 (.A(n_209), .B(n_44), .ZN(p_0[53]));
   XNOR2_X1 i_72 (.A(n_213), .B(n_40), .ZN(p_0[54]));
   XNOR2_X1 i_74 (.A(n_217), .B(n_36), .ZN(p_0[55]));
   XNOR2_X1 i_75 (.A(n_221), .B(n_32), .ZN(p_0[56]));
   XNOR2_X1 i_76 (.A(n_225), .B(n_28), .ZN(p_0[57]));
   XNOR2_X1 i_78 (.A(n_229), .B(n_24), .ZN(p_0[58]));
   XNOR2_X1 i_79 (.A(n_233), .B(n_20), .ZN(p_0[59]));
   XNOR2_X1 i_80 (.A(n_237), .B(n_16), .ZN(p_0[60]));
   XNOR2_X1 i_82 (.A(n_241), .B(n_12), .ZN(p_0[61]));
   XNOR2_X1 i_83 (.A(n_245), .B(n_8), .ZN(p_0[62]));
   XOR2_X1 i_84 (.A(n_4), .B(n_3), .Z(p_0[63]));
   XNOR2_X1 i_86 (.A(partialProd[63]), .B(Acc[63]), .ZN(n_3));
   AOI21_X1 i_87 (.A(n_246), .B1(n_245), .B2(n_7), .ZN(n_4));
   INV_X1 i_88 (.A(n_8), .ZN(n_7));
   AOI21_X1 i_90 (.A(n_242), .B1(n_241), .B2(n_11), .ZN(n_8));
   INV_X1 i_91 (.A(n_12), .ZN(n_11));
   AOI21_X1 i_92 (.A(n_238), .B1(n_237), .B2(n_15), .ZN(n_12));
   INV_X1 i_94 (.A(n_16), .ZN(n_15));
   AOI21_X1 i_95 (.A(n_234), .B1(n_233), .B2(n_19), .ZN(n_16));
   INV_X1 i_96 (.A(n_20), .ZN(n_19));
   AOI21_X1 i_98 (.A(n_230), .B1(n_229), .B2(n_23), .ZN(n_20));
   INV_X1 i_99 (.A(n_24), .ZN(n_23));
   AOI21_X1 i_100 (.A(n_226), .B1(n_225), .B2(n_27), .ZN(n_24));
   INV_X1 i_102 (.A(n_28), .ZN(n_27));
   AOI21_X1 i_103 (.A(n_222), .B1(n_221), .B2(n_31), .ZN(n_28));
   INV_X1 i_104 (.A(n_32), .ZN(n_31));
   AOI21_X1 i_106 (.A(n_218), .B1(n_217), .B2(n_35), .ZN(n_32));
   INV_X1 i_107 (.A(n_36), .ZN(n_35));
   AOI21_X1 i_108 (.A(n_214), .B1(n_213), .B2(n_39), .ZN(n_36));
   INV_X1 i_110 (.A(n_40), .ZN(n_39));
   AOI21_X1 i_111 (.A(n_210), .B1(n_209), .B2(n_43), .ZN(n_40));
   INV_X1 i_112 (.A(n_44), .ZN(n_43));
   AOI21_X1 i_114 (.A(n_206), .B1(n_205), .B2(n_47), .ZN(n_44));
   INV_X1 i_115 (.A(n_48), .ZN(n_47));
   AOI21_X1 i_116 (.A(n_202), .B1(n_201), .B2(n_51), .ZN(n_48));
   INV_X1 i_118 (.A(n_52), .ZN(n_51));
   AOI21_X1 i_119 (.A(n_198), .B1(n_197), .B2(n_55), .ZN(n_52));
   INV_X1 i_120 (.A(n_56), .ZN(n_55));
   AOI21_X1 i_122 (.A(n_194), .B1(n_193), .B2(n_59), .ZN(n_56));
   INV_X1 i_123 (.A(n_60), .ZN(n_59));
   AOI21_X1 i_124 (.A(n_190), .B1(n_189), .B2(n_63), .ZN(n_60));
   INV_X1 i_126 (.A(n_64), .ZN(n_63));
   AOI21_X1 i_127 (.A(n_186), .B1(n_185), .B2(n_67), .ZN(n_64));
   INV_X1 i_128 (.A(n_68), .ZN(n_67));
   AOI21_X1 i_130 (.A(n_182), .B1(n_181), .B2(n_71), .ZN(n_68));
   INV_X1 i_131 (.A(n_72), .ZN(n_71));
   AOI21_X1 i_132 (.A(n_178), .B1(n_177), .B2(n_75), .ZN(n_72));
   INV_X1 i_134 (.A(n_76), .ZN(n_75));
   AOI21_X1 i_135 (.A(n_174), .B1(n_173), .B2(n_79), .ZN(n_76));
   INV_X1 i_136 (.A(n_80), .ZN(n_79));
   AOI21_X1 i_138 (.A(n_170), .B1(n_169), .B2(n_83), .ZN(n_80));
   INV_X1 i_139 (.A(n_84), .ZN(n_83));
   AOI21_X1 i_140 (.A(n_166), .B1(n_165), .B2(n_87), .ZN(n_84));
   INV_X1 i_142 (.A(n_88), .ZN(n_87));
   AOI21_X1 i_143 (.A(n_162), .B1(n_161), .B2(n_91), .ZN(n_88));
   INV_X1 i_144 (.A(n_92), .ZN(n_91));
   AOI21_X1 i_146 (.A(n_158), .B1(n_157), .B2(n_95), .ZN(n_92));
   INV_X1 i_147 (.A(n_96), .ZN(n_95));
   AOI21_X1 i_148 (.A(n_154), .B1(n_153), .B2(n_99), .ZN(n_96));
   INV_X1 i_150 (.A(n_100), .ZN(n_99));
   AOI21_X1 i_151 (.A(n_150), .B1(n_149), .B2(n_103), .ZN(n_100));
   INV_X1 i_152 (.A(n_104), .ZN(n_103));
   AOI21_X1 i_154 (.A(n_146), .B1(n_145), .B2(n_107), .ZN(n_104));
   INV_X1 i_155 (.A(n_108), .ZN(n_107));
   AOI21_X1 i_156 (.A(n_142), .B1(n_141), .B2(n_111), .ZN(n_108));
   INV_X1 i_158 (.A(n_112), .ZN(n_111));
   AOI21_X1 i_159 (.A(n_138), .B1(n_137), .B2(n_115), .ZN(n_112));
   INV_X1 i_160 (.A(n_116), .ZN(n_115));
   AOI21_X1 i_162 (.A(n_134), .B1(n_133), .B2(n_119), .ZN(n_116));
   INV_X1 i_163 (.A(n_120), .ZN(n_119));
   AOI21_X1 i_164 (.A(n_130), .B1(n_129), .B2(n_123), .ZN(n_120));
   INV_X1 i_166 (.A(n_124), .ZN(n_123));
   AOI21_X1 i_167 (.A(n_126), .B1(n_125), .B2(n_127), .ZN(n_124));
   INV_X1 i_168 (.A(n_128), .ZN(n_127));
   AOI21_X1 i_170 (.A(n_122), .B1(n_121), .B2(n_131), .ZN(n_128));
   INV_X1 i_171 (.A(n_132), .ZN(n_131));
   AOI21_X1 i_172 (.A(n_118), .B1(n_117), .B2(n_135), .ZN(n_132));
   INV_X1 i_174 (.A(n_136), .ZN(n_135));
   AOI21_X1 i_175 (.A(n_114), .B1(n_113), .B2(n_139), .ZN(n_136));
   INV_X1 i_176 (.A(n_140), .ZN(n_139));
   AOI21_X1 i_178 (.A(n_110), .B1(n_109), .B2(n_143), .ZN(n_140));
   INV_X1 i_179 (.A(n_144), .ZN(n_143));
   AOI21_X1 i_180 (.A(n_106), .B1(n_105), .B2(n_147), .ZN(n_144));
   INV_X1 i_182 (.A(n_148), .ZN(n_147));
   AOI21_X1 i_183 (.A(n_102), .B1(n_101), .B2(n_151), .ZN(n_148));
   INV_X1 i_184 (.A(n_152), .ZN(n_151));
   AOI21_X1 i_186 (.A(n_98), .B1(n_97), .B2(n_155), .ZN(n_152));
   INV_X1 i_187 (.A(n_156), .ZN(n_155));
   AOI21_X1 i_188 (.A(n_94), .B1(n_93), .B2(n_159), .ZN(n_156));
   INV_X1 i_190 (.A(n_160), .ZN(n_159));
   AOI21_X1 i_191 (.A(n_90), .B1(n_89), .B2(n_163), .ZN(n_160));
   INV_X1 i_192 (.A(n_164), .ZN(n_163));
   AOI21_X1 i_194 (.A(n_86), .B1(n_85), .B2(n_167), .ZN(n_164));
   INV_X1 i_195 (.A(n_168), .ZN(n_167));
   AOI21_X1 i_196 (.A(n_82), .B1(n_81), .B2(n_171), .ZN(n_168));
   INV_X1 i_198 (.A(n_172), .ZN(n_171));
   AOI21_X1 i_199 (.A(n_78), .B1(n_77), .B2(n_175), .ZN(n_172));
   INV_X1 i_200 (.A(n_176), .ZN(n_175));
   AOI21_X1 i_202 (.A(n_74), .B1(n_73), .B2(n_179), .ZN(n_176));
   INV_X1 i_203 (.A(n_180), .ZN(n_179));
   AOI21_X1 i_204 (.A(n_70), .B1(n_69), .B2(n_183), .ZN(n_180));
   INV_X1 i_206 (.A(n_184), .ZN(n_183));
   AOI21_X1 i_207 (.A(n_66), .B1(n_65), .B2(n_187), .ZN(n_184));
   INV_X1 i_208 (.A(n_188), .ZN(n_187));
   AOI21_X1 i_210 (.A(n_62), .B1(n_61), .B2(n_191), .ZN(n_188));
   INV_X1 i_211 (.A(n_192), .ZN(n_191));
   AOI21_X1 i_212 (.A(n_58), .B1(n_57), .B2(n_195), .ZN(n_192));
   INV_X1 i_214 (.A(n_196), .ZN(n_195));
   AOI21_X1 i_215 (.A(n_54), .B1(n_53), .B2(n_199), .ZN(n_196));
   INV_X1 i_216 (.A(n_200), .ZN(n_199));
   AOI21_X1 i_218 (.A(n_50), .B1(n_49), .B2(n_203), .ZN(n_200));
   INV_X1 i_219 (.A(n_204), .ZN(n_203));
   AOI21_X1 i_220 (.A(n_46), .B1(n_45), .B2(n_207), .ZN(n_204));
   INV_X1 i_222 (.A(n_208), .ZN(n_207));
   AOI21_X1 i_223 (.A(n_42), .B1(n_41), .B2(n_211), .ZN(n_208));
   INV_X1 i_224 (.A(n_212), .ZN(n_211));
   AOI21_X1 i_226 (.A(n_38), .B1(n_37), .B2(n_215), .ZN(n_212));
   INV_X1 i_227 (.A(n_216), .ZN(n_215));
   AOI21_X1 i_228 (.A(n_34), .B1(n_33), .B2(n_219), .ZN(n_216));
   INV_X1 i_230 (.A(n_220), .ZN(n_219));
   AOI21_X1 i_231 (.A(n_30), .B1(n_29), .B2(n_223), .ZN(n_220));
   INV_X1 i_232 (.A(n_224), .ZN(n_223));
   AOI21_X1 i_234 (.A(n_26), .B1(n_25), .B2(n_227), .ZN(n_224));
   INV_X1 i_235 (.A(n_228), .ZN(n_227));
   AOI21_X1 i_236 (.A(n_22), .B1(n_21), .B2(n_231), .ZN(n_228));
   INV_X1 i_238 (.A(n_232), .ZN(n_231));
   AOI21_X1 i_239 (.A(n_18), .B1(n_17), .B2(n_235), .ZN(n_232));
   INV_X1 i_240 (.A(n_236), .ZN(n_235));
   AOI21_X1 i_242 (.A(n_14), .B1(n_13), .B2(n_239), .ZN(n_236));
   INV_X1 i_243 (.A(n_240), .ZN(n_239));
   AOI21_X1 i_244 (.A(n_10), .B1(n_9), .B2(n_243), .ZN(n_240));
   INV_X1 i_246 (.A(n_244), .ZN(n_243));
   AOI21_X1 i_247 (.A(n_6), .B1(n_5), .B2(n_247), .ZN(n_244));
   INV_X1 i_248 (.A(n_248), .ZN(n_247));
   AOI21_X1 i_249 (.A(n_2), .B1(n_0), .B2(n_1), .ZN(n_248));
endmodule

module Booth(inputA, inputB, result, clk, reset, en, start);
   input [31:0]inputA;
   input [31:0]inputB;
   output [63:0]result;
   input clk;
   input reset;
   input en;
   input start;

   wire [31:0]B_reg;
   wire [31:0]A_reg;
   wire n_0_0;
   wire [63:0]out_reg;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_0_4;
   wire n_0_0_0;
   wire n_0_0_5;
   wire n_0_0_1;
   wire n_0_0_6;
   wire n_0_0_2;
   wire n_0_0_7;
   wire n_0_0_3;
   wire n_0_0_8;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire [63:0]partialProd;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_443;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_0_481;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_484;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_491;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_0_494;
   wire n_0_0_495;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_502;
   wire n_0_0_503;
   wire n_0_0_504;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_0_512;
   wire n_0_0_513;
   wire n_0_0_514;
   wire n_0_0_515;
   wire n_0_0_516;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_0_526;
   wire n_0_0_527;
   wire n_0_0_528;
   wire n_0_0_529;
   wire n_0_0_530;
   wire n_0_0_531;
   wire n_0_0_532;
   wire n_0_0_533;
   wire n_0_0_534;
   wire n_0_0_535;
   wire n_0_0_536;
   wire n_0_0_537;
   wire n_0_0_538;
   wire n_0_0_539;
   wire n_0_0_540;
   wire n_0_0_541;
   wire n_0_0_542;
   wire n_0_0_543;
   wire n_0_0_544;
   wire n_0_0_545;
   wire n_0_0_546;
   wire n_0_0_547;
   wire n_0_0_548;
   wire n_0_0_549;
   wire n_0_0_550;
   wire n_0_0_551;
   wire n_0_0_552;
   wire n_0_0_553;
   wire n_0_0_554;
   wire n_0_0_555;
   wire n_0_0_556;
   wire n_0_0_557;
   wire n_0_0_558;
   wire n_0_0_559;
   wire n_0_0_560;
   wire n_0_0_561;
   wire n_0_0_562;
   wire n_0_0_563;
   wire n_0_0_564;
   wire n_0_0_565;
   wire n_0_0_566;
   wire n_0_0_567;
   wire n_0_0_568;
   wire n_0_0_569;
   wire n_0_0_570;
   wire n_0_0_571;
   wire n_0_0_572;
   wire n_0_0_573;
   wire n_0_0_574;
   wire n_0_0_575;
   wire n_0_0_576;
   wire n_0_0_577;
   wire n_0_0_578;
   wire n_0_0_579;
   wire n_0_0_580;
   wire n_0_0_581;
   wire n_0_0_582;
   wire n_0_0_583;
   wire n_0_0_584;
   wire n_0_0_585;
   wire n_0_0_586;
   wire n_0_0_587;
   wire n_0_0_588;
   wire n_0_0_589;
   wire n_0_0_590;
   wire n_0_0_591;
   wire n_0_0_592;
   wire n_0_0_593;
   wire n_0_0_594;
   wire n_0_0_595;
   wire n_0_0_596;
   wire n_0_0_597;
   wire n_0_0_598;
   wire n_0_0_599;
   wire n_0_0_600;
   wire n_0_0_601;
   wire n_0_0_602;
   wire n_0_0_603;
   wire n_0_0_604;
   wire n_0_0_605;
   wire n_0_0_606;
   wire n_0_0_607;
   wire n_0_0_608;
   wire n_0_0_609;
   wire n_0_0_610;
   wire n_0_0_611;
   wire n_0_0_612;
   wire n_0_0_613;
   wire n_0_0_614;
   wire n_0_0_615;
   wire n_0_0_616;
   wire n_0_0_617;
   wire n_0_0_618;
   wire n_0_0_619;
   wire n_0_0_620;
   wire n_0_0_621;
   wire n_0_0_622;
   wire n_0_0_623;
   wire n_0_0_624;
   wire n_0_0_625;
   wire n_0_0_626;
   wire n_0_0_627;
   wire n_0_0_628;
   wire n_0_0_629;
   wire n_0_0_630;
   wire n_0_0_631;
   wire n_0_0_632;
   wire n_0_0_633;
   wire n_0_0_634;
   wire n_0_0_635;
   wire n_0_0_636;
   wire n_0_0_637;
   wire n_0_0_638;
   wire n_0_0_639;
   wire n_0_0_640;
   wire n_0_0_641;
   wire n_0_0_642;
   wire n_0_0_643;
   wire n_0_0_644;
   wire n_0_0_645;
   wire n_0_0_646;
   wire n_0_0_647;
   wire n_0_0_648;
   wire n_0_0_649;
   wire n_0_0_650;
   wire n_0_0_651;
   wire n_0_0_652;
   wire n_0_0_653;
   wire n_0_0_654;
   wire n_0_0_655;
   wire n_0_0_656;
   wire n_0_0_657;
   wire n_0_0_658;
   wire n_0_0_659;
   wire n_0_0_660;
   wire n_0_0_661;
   wire n_0_0_662;
   wire n_0_0_663;
   wire n_0_0_664;
   wire n_0_0_665;
   wire n_0_0_666;
   wire n_0_0_667;
   wire n_0_0_668;
   wire n_0_0_669;
   wire n_0_0_670;
   wire n_0_0_671;
   wire n_0_0_672;
   wire n_0_0_673;
   wire n_0_0_674;
   wire n_0_0_675;
   wire n_0_0_676;
   wire n_0_0_677;
   wire n_0_0_678;
   wire n_0_0_679;
   wire n_0_0_680;
   wire n_0_0_681;
   wire n_0_0_682;
   wire n_0_0_683;
   wire n_0_0_684;
   wire n_0_0_685;
   wire n_0_0_686;
   wire n_0_0_687;
   wire n_0_0_688;
   wire n_0_0_689;
   wire n_0_0_690;
   wire n_0_0_691;
   wire n_0_0_692;
   wire n_0_0_693;
   wire n_0_0_694;
   wire n_0_0_695;
   wire n_0_0_696;
   wire n_0_0_697;
   wire n_0_0_698;
   wire n_0_0_699;
   wire n_0_0_700;
   wire n_0_0_701;
   wire n_0_0_702;
   wire n_0_0_703;
   wire n_0_0_704;
   wire n_0_0_705;
   wire n_0_0_706;
   wire n_0_0_707;
   wire n_0_0_708;
   wire n_0_0_709;
   wire n_0_0_710;
   wire n_0_0_711;
   wire n_0_0_712;
   wire n_0_0_713;
   wire n_0_0_714;
   wire n_0_0_715;
   wire n_0_0_716;
   wire n_0_0_717;
   wire n_0_0_718;
   wire n_0_0_719;
   wire n_0_0_720;
   wire n_0_0_721;
   wire n_0_0_722;
   wire n_0_0_723;
   wire n_0_0_724;
   wire n_0_0_725;
   wire n_0_0_726;
   wire n_0_0_727;
   wire n_0_0_728;
   wire n_0_0_729;
   wire n_0_0_730;
   wire n_0_0_731;
   wire n_0_0_732;
   wire n_0_0_733;
   wire n_0_0_734;
   wire n_0_0_735;
   wire n_0_0_736;
   wire n_0_0_737;
   wire n_0_0_738;
   wire n_0_0_739;
   wire n_0_0_740;
   wire n_0_0_741;
   wire n_0_0_742;
   wire n_0_0_743;
   wire n_0_0_744;
   wire n_0_0_745;
   wire n_0_0_746;
   wire n_0_0_747;
   wire n_0_0_748;
   wire n_0_0_749;
   wire n_0_0_750;
   wire n_0_0_751;
   wire n_0_0_752;
   wire n_0_0_753;
   wire n_0_0_754;
   wire n_0_0_755;
   wire n_0_0_756;
   wire n_0_0_757;
   wire n_0_0_758;
   wire n_0_0_759;
   wire n_0_0_760;
   wire n_0_0_761;
   wire n_0_0_762;
   wire n_0_0_763;
   wire n_0_0_764;
   wire n_0_0_765;
   wire n_0_0_766;
   wire n_0_0_767;
   wire n_0_0_768;
   wire n_0_0_769;
   wire n_0_0_770;
   wire n_0_0_771;
   wire n_0_0_772;
   wire n_0_0_773;
   wire n_0_0_774;
   wire n_0_0_775;
   wire n_0_0_776;
   wire n_0_0_777;
   wire n_0_0_778;
   wire n_0_0_779;
   wire n_0_0_780;
   wire n_0_0_781;
   wire n_0_0_782;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_0_783;
   wire n_0_167;
   wire n_0_162;
   wire n_0_169;
   wire n_0_168;
   wire [63:0]Acc;
   wire [63:0]extended_M_mul_neg_one;
   wire [5:0]i;
   wire [63:0]extended_M;
   wire [32:0]Q;
   wire n_0_1;
   wire n_0_33;

   registerNbits__0_16 regB (.clk(clk), .reset(reset), .en(en), .inp(inputB), 
      .out(B_reg));
   registerNbits regA (.clk(clk), .reset(reset), .en(en), .inp(inputA), .out(
      A_reg));
   registerNbits__parameterized0 regOut (.clk(clk), .reset(reset), .en(en), 
      .inp(out_reg), .out(result));
   CLKGATETST_X1 clk_gate_out_reg_reg (.CK(clk), .E(n_0_169), .SE(1'b0), 
      .GCK(n_0_0));
   DFF_X1 \out_reg_reg[63]  (.D(Acc[63]), .CK(n_0_0), .Q(out_reg[63]), .QN());
   DFF_X1 \out_reg_reg[62]  (.D(Acc[62]), .CK(n_0_0), .Q(out_reg[62]), .QN());
   DFF_X1 \out_reg_reg[61]  (.D(Acc[61]), .CK(n_0_0), .Q(out_reg[61]), .QN());
   DFF_X1 \out_reg_reg[60]  (.D(Acc[60]), .CK(n_0_0), .Q(out_reg[60]), .QN());
   DFF_X1 \out_reg_reg[59]  (.D(Acc[59]), .CK(n_0_0), .Q(out_reg[59]), .QN());
   DFF_X1 \out_reg_reg[58]  (.D(Acc[58]), .CK(n_0_0), .Q(out_reg[58]), .QN());
   DFF_X1 \out_reg_reg[57]  (.D(Acc[57]), .CK(n_0_0), .Q(out_reg[57]), .QN());
   DFF_X1 \out_reg_reg[56]  (.D(Acc[56]), .CK(n_0_0), .Q(out_reg[56]), .QN());
   DFF_X1 \out_reg_reg[55]  (.D(Acc[55]), .CK(n_0_0), .Q(out_reg[55]), .QN());
   DFF_X1 \out_reg_reg[54]  (.D(Acc[54]), .CK(n_0_0), .Q(out_reg[54]), .QN());
   DFF_X1 \out_reg_reg[53]  (.D(Acc[53]), .CK(n_0_0), .Q(out_reg[53]), .QN());
   DFF_X1 \out_reg_reg[52]  (.D(Acc[52]), .CK(n_0_0), .Q(out_reg[52]), .QN());
   DFF_X1 \out_reg_reg[51]  (.D(Acc[51]), .CK(n_0_0), .Q(out_reg[51]), .QN());
   DFF_X1 \out_reg_reg[50]  (.D(Acc[50]), .CK(n_0_0), .Q(out_reg[50]), .QN());
   DFF_X1 \out_reg_reg[49]  (.D(Acc[49]), .CK(n_0_0), .Q(out_reg[49]), .QN());
   DFF_X1 \out_reg_reg[48]  (.D(Acc[48]), .CK(n_0_0), .Q(out_reg[48]), .QN());
   DFF_X1 \out_reg_reg[47]  (.D(Acc[47]), .CK(n_0_0), .Q(out_reg[47]), .QN());
   DFF_X1 \out_reg_reg[46]  (.D(Acc[46]), .CK(n_0_0), .Q(out_reg[46]), .QN());
   DFF_X1 \out_reg_reg[45]  (.D(Acc[45]), .CK(n_0_0), .Q(out_reg[45]), .QN());
   DFF_X1 \out_reg_reg[44]  (.D(Acc[44]), .CK(n_0_0), .Q(out_reg[44]), .QN());
   DFF_X1 \out_reg_reg[43]  (.D(Acc[43]), .CK(n_0_0), .Q(out_reg[43]), .QN());
   DFF_X1 \out_reg_reg[42]  (.D(Acc[42]), .CK(n_0_0), .Q(out_reg[42]), .QN());
   DFF_X1 \out_reg_reg[41]  (.D(Acc[41]), .CK(n_0_0), .Q(out_reg[41]), .QN());
   DFF_X1 \out_reg_reg[40]  (.D(Acc[40]), .CK(n_0_0), .Q(out_reg[40]), .QN());
   DFF_X1 \out_reg_reg[39]  (.D(Acc[39]), .CK(n_0_0), .Q(out_reg[39]), .QN());
   DFF_X1 \out_reg_reg[38]  (.D(Acc[38]), .CK(n_0_0), .Q(out_reg[38]), .QN());
   DFF_X1 \out_reg_reg[37]  (.D(Acc[37]), .CK(n_0_0), .Q(out_reg[37]), .QN());
   DFF_X1 \out_reg_reg[36]  (.D(Acc[36]), .CK(n_0_0), .Q(out_reg[36]), .QN());
   DFF_X1 \out_reg_reg[35]  (.D(Acc[35]), .CK(n_0_0), .Q(out_reg[35]), .QN());
   DFF_X1 \out_reg_reg[34]  (.D(Acc[34]), .CK(n_0_0), .Q(out_reg[34]), .QN());
   DFF_X1 \out_reg_reg[33]  (.D(Acc[33]), .CK(n_0_0), .Q(out_reg[33]), .QN());
   DFF_X1 \out_reg_reg[32]  (.D(Acc[32]), .CK(n_0_0), .Q(out_reg[32]), .QN());
   DFF_X1 \out_reg_reg[31]  (.D(Acc[31]), .CK(n_0_0), .Q(out_reg[31]), .QN());
   DFF_X1 \out_reg_reg[30]  (.D(Acc[30]), .CK(n_0_0), .Q(out_reg[30]), .QN());
   DFF_X1 \out_reg_reg[29]  (.D(Acc[29]), .CK(n_0_0), .Q(out_reg[29]), .QN());
   DFF_X1 \out_reg_reg[28]  (.D(Acc[28]), .CK(n_0_0), .Q(out_reg[28]), .QN());
   DFF_X1 \out_reg_reg[27]  (.D(Acc[27]), .CK(n_0_0), .Q(out_reg[27]), .QN());
   DFF_X1 \out_reg_reg[26]  (.D(Acc[26]), .CK(n_0_0), .Q(out_reg[26]), .QN());
   DFF_X1 \out_reg_reg[25]  (.D(Acc[25]), .CK(n_0_0), .Q(out_reg[25]), .QN());
   DFF_X1 \out_reg_reg[24]  (.D(Acc[24]), .CK(n_0_0), .Q(out_reg[24]), .QN());
   DFF_X1 \out_reg_reg[23]  (.D(Acc[23]), .CK(n_0_0), .Q(out_reg[23]), .QN());
   DFF_X1 \out_reg_reg[22]  (.D(Acc[22]), .CK(n_0_0), .Q(out_reg[22]), .QN());
   DFF_X1 \out_reg_reg[21]  (.D(Acc[21]), .CK(n_0_0), .Q(out_reg[21]), .QN());
   DFF_X1 \out_reg_reg[20]  (.D(Acc[20]), .CK(n_0_0), .Q(out_reg[20]), .QN());
   DFF_X1 \out_reg_reg[19]  (.D(Acc[19]), .CK(n_0_0), .Q(out_reg[19]), .QN());
   DFF_X1 \out_reg_reg[18]  (.D(Acc[18]), .CK(n_0_0), .Q(out_reg[18]), .QN());
   DFF_X1 \out_reg_reg[17]  (.D(Acc[17]), .CK(n_0_0), .Q(out_reg[17]), .QN());
   DFF_X1 \out_reg_reg[16]  (.D(Acc[16]), .CK(n_0_0), .Q(out_reg[16]), .QN());
   DFF_X1 \out_reg_reg[15]  (.D(Acc[15]), .CK(n_0_0), .Q(out_reg[15]), .QN());
   DFF_X1 \out_reg_reg[14]  (.D(Acc[14]), .CK(n_0_0), .Q(out_reg[14]), .QN());
   DFF_X1 \out_reg_reg[13]  (.D(Acc[13]), .CK(n_0_0), .Q(out_reg[13]), .QN());
   DFF_X1 \out_reg_reg[12]  (.D(Acc[12]), .CK(n_0_0), .Q(out_reg[12]), .QN());
   DFF_X1 \out_reg_reg[11]  (.D(Acc[11]), .CK(n_0_0), .Q(out_reg[11]), .QN());
   DFF_X1 \out_reg_reg[10]  (.D(Acc[10]), .CK(n_0_0), .Q(out_reg[10]), .QN());
   DFF_X1 \out_reg_reg[9]  (.D(Acc[9]), .CK(n_0_0), .Q(out_reg[9]), .QN());
   DFF_X1 \out_reg_reg[8]  (.D(Acc[8]), .CK(n_0_0), .Q(out_reg[8]), .QN());
   DFF_X1 \out_reg_reg[7]  (.D(Acc[7]), .CK(n_0_0), .Q(out_reg[7]), .QN());
   DFF_X1 \out_reg_reg[6]  (.D(Acc[6]), .CK(n_0_0), .Q(out_reg[6]), .QN());
   DFF_X1 \out_reg_reg[5]  (.D(Acc[5]), .CK(n_0_0), .Q(out_reg[5]), .QN());
   DFF_X1 \out_reg_reg[4]  (.D(Acc[4]), .CK(n_0_0), .Q(out_reg[4]), .QN());
   DFF_X1 \out_reg_reg[3]  (.D(Acc[3]), .CK(n_0_0), .Q(out_reg[3]), .QN());
   DFF_X1 \out_reg_reg[2]  (.D(Acc[2]), .CK(n_0_0), .Q(out_reg[2]), .QN());
   DFF_X1 \out_reg_reg[1]  (.D(Acc[1]), .CK(n_0_0), .Q(out_reg[1]), .QN());
   DFF_X1 \out_reg_reg[0]  (.D(Acc[0]), .CK(n_0_0), .Q(out_reg[0]), .QN());
   datapath i_0_1 (.p_0({n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
      n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
      n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, uc_0}), .A_reg(A_reg));
   datapath__0_12 i_0_10 (.partialProd(partialProd), .Acc(Acc), .p_0({n_0_97, 
      n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, 
      n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, 
      n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, 
      n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, 
      n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, 
      n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, 
      n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34}));
   HA_X1 i_0_0_0 (.A(i[1]), .B(i[0]), .CO(n_0_0_0), .S(n_0_0_4));
   HA_X1 i_0_0_1 (.A(i[2]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_5));
   HA_X1 i_0_0_2 (.A(i[3]), .B(n_0_0_1), .CO(n_0_0_2), .S(n_0_0_6));
   HA_X1 i_0_0_3 (.A(i[4]), .B(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_7));
   INV_X1 i_0_0_4 (.A(start), .ZN(n_0_0_8));
   AND2_X1 i_0_0_5 (.A1(n_0_0_8), .A2(n_0_34), .ZN(n_0_98));
   AND2_X1 i_0_0_6 (.A1(n_0_0_8), .A2(n_0_35), .ZN(n_0_99));
   AND2_X1 i_0_0_7 (.A1(n_0_0_8), .A2(n_0_36), .ZN(n_0_100));
   AND2_X1 i_0_0_8 (.A1(n_0_0_8), .A2(n_0_37), .ZN(n_0_101));
   AND2_X1 i_0_0_9 (.A1(n_0_0_8), .A2(n_0_38), .ZN(n_0_102));
   AND2_X1 i_0_0_10 (.A1(n_0_0_8), .A2(n_0_39), .ZN(n_0_103));
   AND2_X1 i_0_0_11 (.A1(n_0_0_8), .A2(n_0_40), .ZN(n_0_104));
   AND2_X1 i_0_0_12 (.A1(n_0_0_8), .A2(n_0_41), .ZN(n_0_105));
   AND2_X1 i_0_0_13 (.A1(n_0_0_8), .A2(n_0_42), .ZN(n_0_106));
   AND2_X1 i_0_0_14 (.A1(n_0_0_8), .A2(n_0_43), .ZN(n_0_107));
   AND2_X1 i_0_0_15 (.A1(n_0_0_8), .A2(n_0_44), .ZN(n_0_108));
   AND2_X1 i_0_0_16 (.A1(n_0_0_8), .A2(n_0_45), .ZN(n_0_109));
   AND2_X1 i_0_0_17 (.A1(n_0_0_8), .A2(n_0_46), .ZN(n_0_110));
   AND2_X1 i_0_0_18 (.A1(n_0_0_8), .A2(n_0_47), .ZN(n_0_111));
   AND2_X1 i_0_0_19 (.A1(n_0_0_8), .A2(n_0_48), .ZN(n_0_112));
   AND2_X1 i_0_0_20 (.A1(n_0_0_8), .A2(n_0_49), .ZN(n_0_113));
   AND2_X1 i_0_0_21 (.A1(n_0_0_8), .A2(n_0_50), .ZN(n_0_114));
   AND2_X1 i_0_0_22 (.A1(n_0_0_8), .A2(n_0_51), .ZN(n_0_115));
   AND2_X1 i_0_0_23 (.A1(n_0_0_8), .A2(n_0_52), .ZN(n_0_116));
   AND2_X1 i_0_0_24 (.A1(n_0_0_8), .A2(n_0_53), .ZN(n_0_117));
   AND2_X1 i_0_0_25 (.A1(n_0_0_8), .A2(n_0_54), .ZN(n_0_118));
   AND2_X1 i_0_0_26 (.A1(n_0_0_8), .A2(n_0_55), .ZN(n_0_119));
   AND2_X1 i_0_0_27 (.A1(n_0_0_8), .A2(n_0_56), .ZN(n_0_120));
   AND2_X1 i_0_0_28 (.A1(n_0_0_8), .A2(n_0_57), .ZN(n_0_121));
   AND2_X1 i_0_0_29 (.A1(n_0_0_8), .A2(n_0_58), .ZN(n_0_122));
   AND2_X1 i_0_0_30 (.A1(n_0_0_8), .A2(n_0_59), .ZN(n_0_123));
   AND2_X1 i_0_0_31 (.A1(n_0_0_8), .A2(n_0_60), .ZN(n_0_124));
   AND2_X1 i_0_0_32 (.A1(n_0_0_8), .A2(n_0_61), .ZN(n_0_125));
   AND2_X1 i_0_0_33 (.A1(n_0_0_8), .A2(n_0_62), .ZN(n_0_126));
   AND2_X1 i_0_0_34 (.A1(n_0_0_8), .A2(n_0_63), .ZN(n_0_127));
   AND2_X1 i_0_0_35 (.A1(n_0_0_8), .A2(n_0_64), .ZN(n_0_128));
   AND2_X1 i_0_0_36 (.A1(n_0_0_8), .A2(n_0_65), .ZN(n_0_129));
   AND2_X1 i_0_0_37 (.A1(n_0_0_8), .A2(n_0_66), .ZN(n_0_130));
   AND2_X1 i_0_0_38 (.A1(n_0_0_8), .A2(n_0_67), .ZN(n_0_131));
   AND2_X1 i_0_0_39 (.A1(n_0_0_8), .A2(n_0_68), .ZN(n_0_132));
   AND2_X1 i_0_0_40 (.A1(n_0_0_8), .A2(n_0_69), .ZN(n_0_133));
   AND2_X1 i_0_0_41 (.A1(n_0_0_8), .A2(n_0_70), .ZN(n_0_134));
   AND2_X1 i_0_0_42 (.A1(n_0_0_8), .A2(n_0_71), .ZN(n_0_135));
   AND2_X1 i_0_0_43 (.A1(n_0_0_8), .A2(n_0_72), .ZN(n_0_136));
   AND2_X1 i_0_0_44 (.A1(n_0_0_8), .A2(n_0_73), .ZN(n_0_137));
   AND2_X1 i_0_0_45 (.A1(n_0_0_8), .A2(n_0_74), .ZN(n_0_138));
   AND2_X1 i_0_0_46 (.A1(n_0_0_8), .A2(n_0_75), .ZN(n_0_139));
   AND2_X1 i_0_0_47 (.A1(n_0_0_8), .A2(n_0_76), .ZN(n_0_140));
   AND2_X1 i_0_0_48 (.A1(n_0_0_8), .A2(n_0_77), .ZN(n_0_141));
   AND2_X1 i_0_0_49 (.A1(n_0_0_8), .A2(n_0_78), .ZN(n_0_142));
   AND2_X1 i_0_0_50 (.A1(n_0_0_8), .A2(n_0_79), .ZN(n_0_143));
   AND2_X1 i_0_0_51 (.A1(n_0_0_8), .A2(n_0_80), .ZN(n_0_144));
   AND2_X1 i_0_0_52 (.A1(n_0_0_8), .A2(n_0_81), .ZN(n_0_145));
   AND2_X1 i_0_0_53 (.A1(n_0_0_8), .A2(n_0_82), .ZN(n_0_146));
   AND2_X1 i_0_0_54 (.A1(n_0_0_8), .A2(n_0_83), .ZN(n_0_147));
   AND2_X1 i_0_0_55 (.A1(n_0_0_8), .A2(n_0_84), .ZN(n_0_148));
   AND2_X1 i_0_0_56 (.A1(n_0_0_8), .A2(n_0_85), .ZN(n_0_149));
   AND2_X1 i_0_0_57 (.A1(n_0_0_8), .A2(n_0_86), .ZN(n_0_150));
   AND2_X1 i_0_0_58 (.A1(n_0_0_8), .A2(n_0_87), .ZN(n_0_151));
   AND2_X1 i_0_0_59 (.A1(n_0_0_8), .A2(n_0_88), .ZN(n_0_152));
   AND2_X1 i_0_0_60 (.A1(n_0_0_8), .A2(n_0_89), .ZN(n_0_153));
   AND2_X1 i_0_0_61 (.A1(n_0_0_8), .A2(n_0_90), .ZN(n_0_154));
   AND2_X1 i_0_0_62 (.A1(n_0_0_8), .A2(n_0_91), .ZN(n_0_155));
   AND2_X1 i_0_0_63 (.A1(n_0_0_8), .A2(n_0_92), .ZN(n_0_156));
   AND2_X1 i_0_0_64 (.A1(n_0_0_8), .A2(n_0_93), .ZN(n_0_157));
   AND2_X1 i_0_0_65 (.A1(n_0_0_8), .A2(n_0_94), .ZN(n_0_158));
   AND2_X1 i_0_0_66 (.A1(n_0_0_8), .A2(n_0_95), .ZN(n_0_159));
   AND2_X1 i_0_0_67 (.A1(n_0_0_8), .A2(n_0_96), .ZN(n_0_160));
   AND2_X1 i_0_0_68 (.A1(n_0_0_8), .A2(n_0_97), .ZN(n_0_161));
   INV_X1 i_0_0_69 (.A(i[3]), .ZN(n_0_0_9));
   INV_X1 i_0_0_70 (.A(i[5]), .ZN(n_0_0_10));
   NAND2_X1 i_0_0_71 (.A1(n_0_0_9), .A2(n_0_0_10), .ZN(n_0_0_11));
   NOR2_X1 i_0_0_72 (.A1(n_0_0_11), .A2(i[4]), .ZN(n_0_0_12));
   NOR2_X1 i_0_0_73 (.A1(i[2]), .A2(i[1]), .ZN(n_0_0_13));
   NAND2_X1 i_0_0_74 (.A1(n_0_0_12), .A2(n_0_0_13), .ZN(n_0_0_14));
   INV_X1 i_0_0_75 (.A(i[0]), .ZN(n_0_0_15));
   NAND2_X1 i_0_0_76 (.A1(n_0_0_15), .A2(extended_M[0]), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_77 (.A1(i[2]), .A2(i[1]), .ZN(n_0_0_17));
   INV_X1 i_0_0_78 (.A(n_0_0_17), .ZN(n_0_0_18));
   INV_X1 i_0_0_79 (.A(i[1]), .ZN(n_0_0_19));
   NAND2_X1 i_0_0_80 (.A1(n_0_0_19), .A2(i[2]), .ZN(n_0_0_20));
   INV_X1 i_0_0_81 (.A(n_0_0_20), .ZN(n_0_0_21));
   AOI222_X1 i_0_0_82 (.A1(n_0_0_18), .A2(Q[24]), .B1(n_0_0_21), .B2(Q[22]), 
      .C1(n_0_0_13), .C2(Q[18]), .ZN(n_0_0_22));
   INV_X1 i_0_0_83 (.A(i[2]), .ZN(n_0_0_23));
   NAND2_X1 i_0_0_84 (.A1(n_0_0_23), .A2(i[1]), .ZN(n_0_0_24));
   INV_X1 i_0_0_85 (.A(n_0_0_24), .ZN(n_0_0_25));
   AOI21_X1 i_0_0_86 (.A(n_0_0_15), .B1(n_0_0_25), .B2(Q[20]), .ZN(n_0_0_26));
   AOI222_X1 i_0_0_87 (.A1(n_0_0_18), .A2(Q[23]), .B1(n_0_0_25), .B2(Q[19]), 
      .C1(n_0_0_13), .C2(Q[17]), .ZN(n_0_0_27));
   AOI21_X1 i_0_0_88 (.A(i[0]), .B1(n_0_0_21), .B2(Q[21]), .ZN(n_0_0_28));
   AOI22_X1 i_0_0_89 (.A1(n_0_0_22), .A2(n_0_0_26), .B1(n_0_0_27), .B2(n_0_0_28), 
      .ZN(n_0_0_29));
   OAI221_X1 i_0_0_90 (.A(n_0_0_21), .B1(Q[29]), .B2(i[0]), .C1(n_0_0_15), 
      .C2(Q[30]), .ZN(n_0_0_30));
   OAI22_X1 i_0_0_91 (.A1(n_0_0_15), .A2(Q[32]), .B1(Q[31]), .B2(i[0]), .ZN(
      n_0_0_31));
   OAI21_X1 i_0_0_92 (.A(n_0_0_30), .B1(n_0_0_17), .B2(n_0_0_31), .ZN(n_0_0_32));
   OAI22_X1 i_0_0_93 (.A1(n_0_0_15), .A2(Q[28]), .B1(Q[27]), .B2(i[0]), .ZN(
      n_0_0_33));
   INV_X1 i_0_0_94 (.A(n_0_0_13), .ZN(n_0_0_34));
   OAI22_X1 i_0_0_95 (.A1(n_0_0_15), .A2(Q[26]), .B1(Q[25]), .B2(i[0]), .ZN(
      n_0_0_35));
   OAI221_X1 i_0_0_96 (.A(i[3]), .B1(n_0_0_33), .B2(n_0_0_24), .C1(n_0_0_34), 
      .C2(n_0_0_35), .ZN(n_0_0_36));
   OAI22_X1 i_0_0_97 (.A1(n_0_0_29), .A2(i[3]), .B1(n_0_0_32), .B2(n_0_0_36), 
      .ZN(n_0_0_37));
   AOI22_X1 i_0_0_98 (.A1(n_0_0_15), .A2(Q[5]), .B1(Q[6]), .B2(i[0]), .ZN(
      n_0_0_38));
   OAI22_X1 i_0_0_99 (.A1(n_0_0_15), .A2(Q[8]), .B1(Q[7]), .B2(i[0]), .ZN(
      n_0_0_39));
   OAI221_X1 i_0_0_100 (.A(n_0_0_9), .B1(n_0_0_38), .B2(n_0_0_20), .C1(n_0_0_39), 
      .C2(n_0_0_17), .ZN(n_0_0_40));
   INV_X1 i_0_0_101 (.A(Q[1]), .ZN(n_0_0_41));
   INV_X1 i_0_0_102 (.A(Q[2]), .ZN(n_0_0_42));
   AOI221_X1 i_0_0_103 (.A(n_0_0_34), .B1(n_0_0_41), .B2(n_0_0_15), .C1(n_0_0_42), 
      .C2(i[0]), .ZN(n_0_0_43));
   INV_X1 i_0_0_104 (.A(Q[4]), .ZN(n_0_0_44));
   INV_X1 i_0_0_105 (.A(Q[3]), .ZN(n_0_0_45));
   AOI221_X1 i_0_0_106 (.A(n_0_0_24), .B1(n_0_0_44), .B2(i[0]), .C1(n_0_0_45), 
      .C2(n_0_0_15), .ZN(n_0_0_46));
   OAI221_X1 i_0_0_107 (.A(n_0_0_21), .B1(Q[13]), .B2(i[0]), .C1(Q[14]), 
      .C2(n_0_0_15), .ZN(n_0_0_47));
   OAI22_X1 i_0_0_108 (.A1(n_0_0_15), .A2(Q[16]), .B1(Q[15]), .B2(i[0]), 
      .ZN(n_0_0_48));
   OAI21_X1 i_0_0_109 (.A(n_0_0_47), .B1(n_0_0_17), .B2(n_0_0_48), .ZN(n_0_0_49));
   AOI22_X1 i_0_0_110 (.A1(n_0_0_15), .A2(Q[9]), .B1(Q[10]), .B2(i[0]), .ZN(
      n_0_0_50));
   AOI22_X1 i_0_0_111 (.A1(n_0_0_15), .A2(Q[11]), .B1(Q[12]), .B2(i[0]), 
      .ZN(n_0_0_51));
   OAI22_X1 i_0_0_112 (.A1(n_0_0_50), .A2(n_0_0_34), .B1(n_0_0_51), .B2(n_0_0_24), 
      .ZN(n_0_0_52));
   OAI33_X1 i_0_0_113 (.A1(n_0_0_40), .A2(n_0_0_43), .A3(n_0_0_46), .B1(n_0_0_49), 
      .B2(n_0_0_9), .B3(n_0_0_52), .ZN(n_0_0_53));
   INV_X1 i_0_0_114 (.A(i[4]), .ZN(n_0_0_54));
   AOI221_X1 i_0_0_115 (.A(i[5]), .B1(n_0_0_37), .B2(i[4]), .C1(n_0_0_53), 
      .C2(n_0_0_54), .ZN(n_0_0_55));
   INV_X1 i_0_0_116 (.A(Q[5]), .ZN(n_0_0_56));
   AOI221_X1 i_0_0_117 (.A(n_0_0_20), .B1(n_0_0_44), .B2(n_0_0_15), .C1(n_0_0_56), 
      .C2(i[0]), .ZN(n_0_0_57));
   NOR2_X1 i_0_0_118 (.A1(n_0_0_34), .A2(n_0_0_41), .ZN(n_0_0_58));
   AOI22_X1 i_0_0_119 (.A1(n_0_0_42), .A2(n_0_0_15), .B1(n_0_0_45), .B2(i[0]), 
      .ZN(n_0_0_59));
   AOI221_X1 i_0_0_120 (.A(n_0_0_57), .B1(i[0]), .B2(n_0_0_58), .C1(n_0_0_25), 
      .C2(n_0_0_59), .ZN(n_0_0_60));
   OAI221_X1 i_0_0_121 (.A(n_0_0_18), .B1(Q[6]), .B2(i[0]), .C1(n_0_0_15), 
      .C2(Q[7]), .ZN(n_0_0_61));
   AOI21_X1 i_0_0_122 (.A(i[4]), .B1(n_0_0_60), .B2(n_0_0_61), .ZN(n_0_0_62));
   INV_X1 i_0_0_123 (.A(Q[16]), .ZN(n_0_0_63));
   INV_X1 i_0_0_124 (.A(Q[17]), .ZN(n_0_0_64));
   AOI22_X1 i_0_0_125 (.A1(n_0_0_63), .A2(n_0_0_15), .B1(n_0_0_64), .B2(i[0]), 
      .ZN(n_0_0_65));
   INV_X1 i_0_0_126 (.A(Q[22]), .ZN(n_0_0_66));
   INV_X1 i_0_0_127 (.A(Q[23]), .ZN(n_0_0_67));
   AOI22_X1 i_0_0_128 (.A1(n_0_0_66), .A2(n_0_0_15), .B1(n_0_0_67), .B2(i[0]), 
      .ZN(n_0_0_68));
   INV_X1 i_0_0_129 (.A(Q[19]), .ZN(n_0_0_69));
   INV_X1 i_0_0_130 (.A(Q[18]), .ZN(n_0_0_70));
   OAI22_X1 i_0_0_131 (.A1(n_0_0_69), .A2(n_0_0_15), .B1(n_0_0_70), .B2(i[0]), 
      .ZN(n_0_0_71));
   OAI222_X1 i_0_0_132 (.A1(n_0_0_65), .A2(n_0_0_34), .B1(n_0_0_68), .B2(
      n_0_0_17), .C1(n_0_0_71), .C2(n_0_0_24), .ZN(n_0_0_72));
   OAI22_X1 i_0_0_133 (.A1(n_0_0_15), .A2(Q[21]), .B1(Q[20]), .B2(i[0]), 
      .ZN(n_0_0_73));
   AOI211_X1 i_0_0_134 (.A(n_0_0_54), .B(n_0_0_72), .C1(n_0_0_21), .C2(n_0_0_73), 
      .ZN(n_0_0_74));
   INV_X1 i_0_0_135 (.A(Q[29]), .ZN(n_0_0_75));
   INV_X1 i_0_0_136 (.A(Q[28]), .ZN(n_0_0_76));
   OAI22_X1 i_0_0_137 (.A1(n_0_0_75), .A2(n_0_0_15), .B1(n_0_0_76), .B2(i[0]), 
      .ZN(n_0_0_77));
   INV_X1 i_0_0_138 (.A(Q[25]), .ZN(n_0_0_78));
   INV_X1 i_0_0_139 (.A(Q[24]), .ZN(n_0_0_79));
   OAI22_X1 i_0_0_140 (.A1(n_0_0_78), .A2(n_0_0_15), .B1(n_0_0_79), .B2(i[0]), 
      .ZN(n_0_0_80));
   OAI221_X1 i_0_0_141 (.A(i[4]), .B1(n_0_0_77), .B2(n_0_0_20), .C1(n_0_0_34), 
      .C2(n_0_0_80), .ZN(n_0_0_81));
   OAI22_X1 i_0_0_142 (.A1(n_0_0_24), .A2(Q[27]), .B1(n_0_0_17), .B2(Q[31]), 
      .ZN(n_0_0_82));
   OAI22_X1 i_0_0_143 (.A1(n_0_0_24), .A2(Q[26]), .B1(n_0_0_17), .B2(Q[30]), 
      .ZN(n_0_0_83));
   AOI221_X1 i_0_0_144 (.A(n_0_0_81), .B1(i[0]), .B2(n_0_0_82), .C1(n_0_0_15), 
      .C2(n_0_0_83), .ZN(n_0_0_84));
   INV_X1 i_0_0_145 (.A(Q[13]), .ZN(n_0_0_85));
   INV_X1 i_0_0_146 (.A(Q[12]), .ZN(n_0_0_86));
   OAI22_X1 i_0_0_147 (.A1(n_0_0_85), .A2(n_0_0_15), .B1(n_0_0_86), .B2(i[0]), 
      .ZN(n_0_0_87));
   INV_X1 i_0_0_148 (.A(Q[9]), .ZN(n_0_0_88));
   INV_X1 i_0_0_149 (.A(Q[8]), .ZN(n_0_0_89));
   OAI22_X1 i_0_0_150 (.A1(n_0_0_88), .A2(n_0_0_15), .B1(n_0_0_89), .B2(i[0]), 
      .ZN(n_0_0_90));
   OAI221_X1 i_0_0_151 (.A(n_0_0_54), .B1(n_0_0_87), .B2(n_0_0_20), .C1(n_0_0_34), 
      .C2(n_0_0_90), .ZN(n_0_0_91));
   OAI22_X1 i_0_0_152 (.A1(n_0_0_15), .A2(Q[15]), .B1(Q[14]), .B2(i[0]), 
      .ZN(n_0_0_92));
   AOI22_X1 i_0_0_153 (.A1(n_0_0_15), .A2(Q[10]), .B1(Q[11]), .B2(i[0]), 
      .ZN(n_0_0_93));
   AOI221_X1 i_0_0_154 (.A(n_0_0_91), .B1(n_0_0_18), .B2(n_0_0_92), .C1(n_0_0_25), 
      .C2(n_0_0_93), .ZN(n_0_0_94));
   OAI33_X1 i_0_0_155 (.A1(n_0_0_62), .A2(n_0_0_74), .A3(i[3]), .B1(n_0_0_84), 
      .B2(n_0_0_94), .B3(n_0_0_9), .ZN(n_0_0_95));
   OR2_X1 i_0_0_156 (.A1(n_0_0_95), .A2(i[5]), .ZN(n_0_0_96));
   NAND2_X1 i_0_0_157 (.A1(n_0_0_9), .A2(i[5]), .ZN(n_0_0_97));
   NOR3_X1 i_0_0_158 (.A1(n_0_0_34), .A2(n_0_0_97), .A3(i[4]), .ZN(n_0_0_98));
   NAND3_X1 i_0_0_159 (.A1(n_0_0_98), .A2(Q[32]), .A3(n_0_0_15), .ZN(n_0_0_99));
   AOI21_X1 i_0_0_160 (.A(n_0_0_55), .B1(n_0_0_96), .B2(n_0_0_99), .ZN(n_0_0_100));
   INV_X1 i_0_0_161 (.A(n_0_0_100), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_162 (.A1(n_0_0_95), .A2(n_0_0_55), .ZN(n_0_0_102));
   AOI211_X1 i_0_0_163 (.A(n_0_0_14), .B(n_0_0_16), .C1(n_0_0_101), .C2(
      n_0_0_102), .ZN(partialProd[0]));
   INV_X1 i_0_0_164 (.A(extended_M[0]), .ZN(n_0_0_103));
   NOR2_X1 i_0_0_165 (.A1(n_0_0_103), .A2(n_0_0_15), .ZN(n_0_0_104));
   AOI21_X1 i_0_0_166 (.A(n_0_0_104), .B1(extended_M[1]), .B2(n_0_0_15), 
      .ZN(n_0_0_105));
   AOI21_X1 i_0_0_167 (.A(n_0_0_104), .B1(extended_M_mul_neg_one[1]), .B2(
      n_0_0_15), .ZN(n_0_0_106));
   OAI33_X1 i_0_0_168 (.A1(n_0_0_101), .A2(n_0_0_14), .A3(n_0_0_105), .B1(
      n_0_0_102), .B2(n_0_0_14), .B3(n_0_0_106), .ZN(partialProd[1]));
   INV_X1 i_0_0_169 (.A(n_0_0_102), .ZN(n_0_0_107));
   INV_X1 i_0_0_170 (.A(extended_M_mul_neg_one[1]), .ZN(n_0_0_108));
   OAI21_X1 i_0_0_171 (.A(i[0]), .B1(n_0_0_14), .B2(n_0_0_108), .ZN(n_0_0_109));
   INV_X1 i_0_0_172 (.A(n_0_0_12), .ZN(n_0_0_110));
   NOR2_X1 i_0_0_173 (.A1(n_0_0_110), .A2(i[2]), .ZN(n_0_0_111));
   NAND2_X1 i_0_0_174 (.A1(n_0_0_111), .A2(i[1]), .ZN(n_0_0_112));
   OR2_X1 i_0_0_175 (.A1(n_0_0_112), .A2(n_0_0_103), .ZN(n_0_0_113));
   INV_X1 i_0_0_176 (.A(extended_M_mul_neg_one[2]), .ZN(n_0_0_114));
   OAI21_X1 i_0_0_177 (.A(n_0_0_113), .B1(n_0_0_114), .B2(n_0_0_14), .ZN(
      n_0_0_115));
   OAI211_X1 i_0_0_178 (.A(n_0_0_107), .B(n_0_0_109), .C1(i[0]), .C2(n_0_0_115), 
      .ZN(n_0_0_116));
   INV_X1 i_0_0_179 (.A(n_0_0_16), .ZN(n_0_0_117));
   INV_X1 i_0_0_180 (.A(extended_M[1]), .ZN(n_0_0_118));
   INV_X1 i_0_0_181 (.A(extended_M[2]), .ZN(n_0_0_119));
   OAI22_X1 i_0_0_182 (.A1(n_0_0_118), .A2(n_0_0_15), .B1(n_0_0_119), .B2(i[0]), 
      .ZN(n_0_0_120));
   OAI221_X1 i_0_0_183 (.A(n_0_0_111), .B1(n_0_0_117), .B2(n_0_0_19), .C1(
      n_0_0_120), .C2(i[1]), .ZN(n_0_0_121));
   OAI21_X1 i_0_0_184 (.A(n_0_0_116), .B1(n_0_0_101), .B2(n_0_0_121), .ZN(
      partialProd[2]));
   OAI211_X1 i_0_0_185 (.A(n_0_0_113), .B(i[0]), .C1(n_0_0_119), .C2(n_0_0_14), 
      .ZN(n_0_0_122));
   INV_X1 i_0_0_186 (.A(n_0_0_111), .ZN(n_0_0_123));
   AOI22_X1 i_0_0_187 (.A1(n_0_0_19), .A2(extended_M[3]), .B1(extended_M[1]), 
      .B2(i[1]), .ZN(n_0_0_124));
   NOR2_X1 i_0_0_188 (.A1(n_0_0_123), .A2(n_0_0_124), .ZN(n_0_0_125));
   OAI211_X1 i_0_0_189 (.A(n_0_0_100), .B(n_0_0_122), .C1(i[0]), .C2(n_0_0_125), 
      .ZN(n_0_0_126));
   AOI22_X1 i_0_0_190 (.A1(n_0_0_19), .A2(extended_M_mul_neg_one[3]), .B1(
      extended_M_mul_neg_one[1]), .B2(i[1]), .ZN(n_0_0_127));
   NOR2_X1 i_0_0_191 (.A1(n_0_0_123), .A2(n_0_0_127), .ZN(n_0_0_128));
   OAI22_X1 i_0_0_192 (.A1(n_0_0_115), .A2(n_0_0_15), .B1(i[0]), .B2(n_0_0_128), 
      .ZN(n_0_0_129));
   OAI21_X1 i_0_0_193 (.A(n_0_0_126), .B1(n_0_0_102), .B2(n_0_0_129), .ZN(
      partialProd[3]));
   NOR2_X1 i_0_0_194 (.A1(n_0_0_110), .A2(n_0_0_23), .ZN(n_0_0_130));
   NAND3_X1 i_0_0_195 (.A1(n_0_0_130), .A2(extended_M[0]), .A3(n_0_0_21), 
      .ZN(n_0_0_131));
   INV_X1 i_0_0_196 (.A(extended_M[4]), .ZN(n_0_0_132));
   OAI221_X1 i_0_0_197 (.A(n_0_0_131), .B1(n_0_0_132), .B2(n_0_0_14), .C1(
      n_0_0_112), .C2(n_0_0_119), .ZN(n_0_0_133));
   OAI221_X1 i_0_0_198 (.A(n_0_0_100), .B1(i[0]), .B2(n_0_0_133), .C1(n_0_0_15), 
      .C2(n_0_0_125), .ZN(n_0_0_134));
   INV_X1 i_0_0_199 (.A(extended_M_mul_neg_one[4]), .ZN(n_0_0_135));
   OAI221_X1 i_0_0_200 (.A(n_0_0_131), .B1(n_0_0_135), .B2(n_0_0_14), .C1(
      n_0_0_112), .C2(n_0_0_114), .ZN(n_0_0_136));
   OAI22_X1 i_0_0_201 (.A1(n_0_0_136), .A2(i[0]), .B1(n_0_0_15), .B2(n_0_0_128), 
      .ZN(n_0_0_137));
   OAI21_X1 i_0_0_202 (.A(n_0_0_134), .B1(n_0_0_102), .B2(n_0_0_137), .ZN(
      partialProd[4]));
   AOI22_X1 i_0_0_203 (.A1(n_0_0_130), .A2(extended_M[1]), .B1(n_0_0_111), 
      .B2(extended_M[5]), .ZN(n_0_0_138));
   INV_X1 i_0_0_204 (.A(extended_M[3]), .ZN(n_0_0_139));
   OAI22_X1 i_0_0_205 (.A1(n_0_0_138), .A2(i[1]), .B1(n_0_0_112), .B2(n_0_0_139), 
      .ZN(n_0_0_140));
   OAI221_X1 i_0_0_206 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_133), .C1(i[0]), 
      .C2(n_0_0_140), .ZN(n_0_0_141));
   AOI22_X1 i_0_0_207 (.A1(n_0_0_130), .A2(extended_M_mul_neg_one[1]), .B1(
      n_0_0_111), .B2(extended_M_mul_neg_one[5]), .ZN(n_0_0_142));
   INV_X1 i_0_0_208 (.A(extended_M_mul_neg_one[3]), .ZN(n_0_0_143));
   OAI22_X1 i_0_0_209 (.A1(n_0_0_142), .A2(i[1]), .B1(n_0_0_112), .B2(n_0_0_143), 
      .ZN(n_0_0_144));
   OAI22_X1 i_0_0_210 (.A1(n_0_0_136), .A2(n_0_0_15), .B1(n_0_0_144), .B2(i[0]), 
      .ZN(n_0_0_145));
   OAI21_X1 i_0_0_211 (.A(n_0_0_141), .B1(n_0_0_102), .B2(n_0_0_145), .ZN(
      partialProd[5]));
   AOI22_X1 i_0_0_212 (.A1(n_0_0_130), .A2(extended_M[2]), .B1(n_0_0_111), 
      .B2(extended_M[6]), .ZN(n_0_0_146));
   AOI21_X1 i_0_0_213 (.A(n_0_0_19), .B1(n_0_0_130), .B2(extended_M[0]), 
      .ZN(n_0_0_147));
   NAND2_X1 i_0_0_214 (.A1(n_0_0_111), .A2(extended_M[4]), .ZN(n_0_0_148));
   AOI22_X1 i_0_0_215 (.A1(n_0_0_146), .A2(n_0_0_19), .B1(n_0_0_147), .B2(
      n_0_0_148), .ZN(n_0_0_149));
   OAI221_X1 i_0_0_216 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_140), .C1(i[0]), 
      .C2(n_0_0_149), .ZN(n_0_0_150));
   AOI22_X1 i_0_0_217 (.A1(n_0_0_130), .A2(extended_M_mul_neg_one[2]), .B1(
      n_0_0_111), .B2(extended_M_mul_neg_one[6]), .ZN(n_0_0_151));
   NAND2_X1 i_0_0_218 (.A1(n_0_0_111), .A2(extended_M_mul_neg_one[4]), .ZN(
      n_0_0_152));
   AOI22_X1 i_0_0_219 (.A1(n_0_0_151), .A2(n_0_0_19), .B1(n_0_0_147), .B2(
      n_0_0_152), .ZN(n_0_0_153));
   OAI22_X1 i_0_0_220 (.A1(n_0_0_144), .A2(n_0_0_15), .B1(n_0_0_153), .B2(i[0]), 
      .ZN(n_0_0_154));
   OAI21_X1 i_0_0_221 (.A(n_0_0_150), .B1(n_0_0_102), .B2(n_0_0_154), .ZN(
      partialProd[6]));
   AOI22_X1 i_0_0_222 (.A1(n_0_0_130), .A2(extended_M[3]), .B1(n_0_0_111), 
      .B2(extended_M[7]), .ZN(n_0_0_155));
   AOI22_X1 i_0_0_223 (.A1(n_0_0_155), .A2(n_0_0_19), .B1(n_0_0_138), .B2(i[1]), 
      .ZN(n_0_0_156));
   OAI221_X1 i_0_0_224 (.A(n_0_0_100), .B1(i[0]), .B2(n_0_0_156), .C1(n_0_0_15), 
      .C2(n_0_0_149), .ZN(n_0_0_157));
   AOI22_X1 i_0_0_225 (.A1(n_0_0_130), .A2(extended_M_mul_neg_one[3]), .B1(
      n_0_0_111), .B2(extended_M_mul_neg_one[7]), .ZN(n_0_0_158));
   AOI22_X1 i_0_0_226 (.A1(n_0_0_158), .A2(n_0_0_19), .B1(n_0_0_142), .B2(i[1]), 
      .ZN(n_0_0_159));
   OAI22_X1 i_0_0_227 (.A1(n_0_0_159), .A2(i[0]), .B1(n_0_0_153), .B2(n_0_0_15), 
      .ZN(n_0_0_160));
   OAI21_X1 i_0_0_228 (.A(n_0_0_157), .B1(n_0_0_102), .B2(n_0_0_160), .ZN(
      partialProd[7]));
   NAND2_X1 i_0_0_229 (.A1(n_0_0_10), .A2(i[3]), .ZN(n_0_0_161));
   NOR2_X1 i_0_0_230 (.A1(n_0_0_161), .A2(i[4]), .ZN(n_0_0_162));
   NAND2_X1 i_0_0_231 (.A1(n_0_0_162), .A2(extended_M[0]), .ZN(n_0_0_163));
   INV_X1 i_0_0_232 (.A(extended_M[8]), .ZN(n_0_0_164));
   OAI21_X1 i_0_0_233 (.A(n_0_0_163), .B1(n_0_0_164), .B2(n_0_0_110), .ZN(
      n_0_0_165));
   AOI22_X1 i_0_0_234 (.A1(n_0_0_165), .A2(n_0_0_23), .B1(extended_M[4]), 
      .B2(n_0_0_130), .ZN(n_0_0_166));
   AOI22_X1 i_0_0_235 (.A1(n_0_0_166), .A2(n_0_0_19), .B1(n_0_0_146), .B2(i[1]), 
      .ZN(n_0_0_167));
   OAI221_X1 i_0_0_236 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_156), .C1(i[0]), 
      .C2(n_0_0_167), .ZN(n_0_0_168));
   INV_X1 i_0_0_237 (.A(extended_M_mul_neg_one[8]), .ZN(n_0_0_169));
   OAI21_X1 i_0_0_238 (.A(n_0_0_163), .B1(n_0_0_169), .B2(n_0_0_110), .ZN(
      n_0_0_170));
   AOI22_X1 i_0_0_239 (.A1(n_0_0_170), .A2(n_0_0_23), .B1(
      extended_M_mul_neg_one[4]), .B2(n_0_0_130), .ZN(n_0_0_171));
   AOI22_X1 i_0_0_240 (.A1(n_0_0_171), .A2(n_0_0_19), .B1(n_0_0_151), .B2(i[1]), 
      .ZN(n_0_0_172));
   OAI22_X1 i_0_0_241 (.A1(n_0_0_172), .A2(i[0]), .B1(n_0_0_159), .B2(n_0_0_15), 
      .ZN(n_0_0_173));
   OAI21_X1 i_0_0_242 (.A(n_0_0_168), .B1(n_0_0_102), .B2(n_0_0_173), .ZN(
      partialProd[8]));
   INV_X1 i_0_0_243 (.A(n_0_0_162), .ZN(n_0_0_174));
   INV_X1 i_0_0_244 (.A(extended_M[9]), .ZN(n_0_0_175));
   OAI22_X1 i_0_0_245 (.A1(n_0_0_174), .A2(n_0_0_118), .B1(n_0_0_110), .B2(
      n_0_0_175), .ZN(n_0_0_176));
   AOI22_X1 i_0_0_246 (.A1(n_0_0_176), .A2(n_0_0_23), .B1(extended_M[5]), 
      .B2(n_0_0_130), .ZN(n_0_0_177));
   OAI22_X1 i_0_0_247 (.A1(n_0_0_177), .A2(i[1]), .B1(n_0_0_155), .B2(n_0_0_19), 
      .ZN(n_0_0_178));
   OAI221_X1 i_0_0_248 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_167), .C1(i[0]), 
      .C2(n_0_0_178), .ZN(n_0_0_179));
   INV_X1 i_0_0_249 (.A(extended_M_mul_neg_one[9]), .ZN(n_0_0_180));
   OAI22_X1 i_0_0_250 (.A1(n_0_0_174), .A2(n_0_0_108), .B1(n_0_0_110), .B2(
      n_0_0_180), .ZN(n_0_0_181));
   AOI22_X1 i_0_0_251 (.A1(n_0_0_181), .A2(n_0_0_23), .B1(
      extended_M_mul_neg_one[5]), .B2(n_0_0_130), .ZN(n_0_0_182));
   OAI22_X1 i_0_0_252 (.A1(n_0_0_182), .A2(i[1]), .B1(n_0_0_158), .B2(n_0_0_19), 
      .ZN(n_0_0_183));
   OAI22_X1 i_0_0_253 (.A1(n_0_0_172), .A2(n_0_0_15), .B1(n_0_0_183), .B2(i[0]), 
      .ZN(n_0_0_184));
   OAI21_X1 i_0_0_254 (.A(n_0_0_179), .B1(n_0_0_102), .B2(n_0_0_184), .ZN(
      partialProd[9]));
   INV_X1 i_0_0_255 (.A(extended_M[10]), .ZN(n_0_0_185));
   OAI22_X1 i_0_0_256 (.A1(n_0_0_174), .A2(n_0_0_119), .B1(n_0_0_110), .B2(
      n_0_0_185), .ZN(n_0_0_186));
   AOI22_X1 i_0_0_257 (.A1(n_0_0_186), .A2(n_0_0_23), .B1(extended_M[6]), 
      .B2(n_0_0_130), .ZN(n_0_0_187));
   OAI22_X1 i_0_0_258 (.A1(i[1]), .A2(n_0_0_187), .B1(n_0_0_166), .B2(n_0_0_19), 
      .ZN(n_0_0_188));
   OAI221_X1 i_0_0_259 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_178), .C1(i[0]), 
      .C2(n_0_0_188), .ZN(n_0_0_189));
   INV_X1 i_0_0_260 (.A(extended_M_mul_neg_one[10]), .ZN(n_0_0_190));
   OAI22_X1 i_0_0_261 (.A1(n_0_0_174), .A2(n_0_0_114), .B1(n_0_0_110), .B2(
      n_0_0_190), .ZN(n_0_0_191));
   AOI22_X1 i_0_0_262 (.A1(n_0_0_191), .A2(n_0_0_23), .B1(
      extended_M_mul_neg_one[6]), .B2(n_0_0_130), .ZN(n_0_0_192));
   OAI22_X1 i_0_0_263 (.A1(i[1]), .A2(n_0_0_192), .B1(n_0_0_171), .B2(n_0_0_19), 
      .ZN(n_0_0_193));
   OAI22_X1 i_0_0_264 (.A1(n_0_0_193), .A2(i[0]), .B1(n_0_0_183), .B2(n_0_0_15), 
      .ZN(n_0_0_194));
   OAI21_X1 i_0_0_265 (.A(n_0_0_189), .B1(n_0_0_102), .B2(n_0_0_194), .ZN(
      partialProd[10]));
   INV_X1 i_0_0_266 (.A(extended_M[11]), .ZN(n_0_0_195));
   OAI22_X1 i_0_0_267 (.A1(n_0_0_174), .A2(n_0_0_139), .B1(n_0_0_110), .B2(
      n_0_0_195), .ZN(n_0_0_196));
   AOI22_X1 i_0_0_268 (.A1(n_0_0_196), .A2(n_0_0_23), .B1(extended_M[7]), 
      .B2(n_0_0_130), .ZN(n_0_0_197));
   OAI22_X1 i_0_0_269 (.A1(n_0_0_177), .A2(n_0_0_19), .B1(n_0_0_197), .B2(i[1]), 
      .ZN(n_0_0_198));
   OAI221_X1 i_0_0_270 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_188), .C1(i[0]), 
      .C2(n_0_0_198), .ZN(n_0_0_199));
   INV_X1 i_0_0_271 (.A(extended_M_mul_neg_one[11]), .ZN(n_0_0_200));
   OAI22_X1 i_0_0_272 (.A1(n_0_0_174), .A2(n_0_0_143), .B1(n_0_0_110), .B2(
      n_0_0_200), .ZN(n_0_0_201));
   AOI22_X1 i_0_0_273 (.A1(n_0_0_201), .A2(n_0_0_23), .B1(
      extended_M_mul_neg_one[7]), .B2(n_0_0_130), .ZN(n_0_0_202));
   OAI22_X1 i_0_0_274 (.A1(n_0_0_182), .A2(n_0_0_19), .B1(n_0_0_202), .B2(i[1]), 
      .ZN(n_0_0_203));
   OAI22_X1 i_0_0_275 (.A1(n_0_0_193), .A2(n_0_0_15), .B1(n_0_0_203), .B2(i[0]), 
      .ZN(n_0_0_204));
   OAI21_X1 i_0_0_276 (.A(n_0_0_199), .B1(n_0_0_102), .B2(n_0_0_204), .ZN(
      partialProd[11]));
   INV_X1 i_0_0_277 (.A(extended_M[12]), .ZN(n_0_0_205));
   OAI22_X1 i_0_0_278 (.A1(n_0_0_174), .A2(n_0_0_132), .B1(n_0_0_110), .B2(
      n_0_0_205), .ZN(n_0_0_206));
   OAI22_X1 i_0_0_279 (.A1(n_0_0_165), .A2(n_0_0_23), .B1(n_0_0_206), .B2(i[2]), 
      .ZN(n_0_0_207));
   AOI22_X1 i_0_0_280 (.A1(n_0_0_207), .A2(n_0_0_19), .B1(n_0_0_187), .B2(i[1]), 
      .ZN(n_0_0_208));
   OAI221_X1 i_0_0_281 (.A(n_0_0_100), .B1(i[0]), .B2(n_0_0_208), .C1(n_0_0_15), 
      .C2(n_0_0_198), .ZN(n_0_0_209));
   INV_X1 i_0_0_282 (.A(extended_M_mul_neg_one[12]), .ZN(n_0_0_210));
   OAI22_X1 i_0_0_283 (.A1(n_0_0_174), .A2(n_0_0_135), .B1(n_0_0_110), .B2(
      n_0_0_210), .ZN(n_0_0_211));
   OAI22_X1 i_0_0_284 (.A1(n_0_0_170), .A2(n_0_0_23), .B1(n_0_0_211), .B2(i[2]), 
      .ZN(n_0_0_212));
   AOI22_X1 i_0_0_285 (.A1(n_0_0_212), .A2(n_0_0_19), .B1(n_0_0_192), .B2(i[1]), 
      .ZN(n_0_0_213));
   OAI22_X1 i_0_0_286 (.A1(n_0_0_213), .A2(i[0]), .B1(n_0_0_203), .B2(n_0_0_15), 
      .ZN(n_0_0_214));
   OAI21_X1 i_0_0_287 (.A(n_0_0_209), .B1(n_0_0_102), .B2(n_0_0_214), .ZN(
      partialProd[12]));
   INV_X1 i_0_0_288 (.A(extended_M[5]), .ZN(n_0_0_215));
   INV_X1 i_0_0_289 (.A(extended_M[13]), .ZN(n_0_0_216));
   OAI22_X1 i_0_0_290 (.A1(n_0_0_174), .A2(n_0_0_215), .B1(n_0_0_110), .B2(
      n_0_0_216), .ZN(n_0_0_217));
   OAI22_X1 i_0_0_291 (.A1(n_0_0_217), .A2(i[2]), .B1(n_0_0_176), .B2(n_0_0_23), 
      .ZN(n_0_0_218));
   AOI22_X1 i_0_0_292 (.A1(n_0_0_218), .A2(n_0_0_19), .B1(n_0_0_197), .B2(i[1]), 
      .ZN(n_0_0_219));
   OAI221_X1 i_0_0_293 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_208), .C1(i[0]), 
      .C2(n_0_0_219), .ZN(n_0_0_220));
   INV_X1 i_0_0_294 (.A(extended_M_mul_neg_one[5]), .ZN(n_0_0_221));
   INV_X1 i_0_0_295 (.A(extended_M_mul_neg_one[13]), .ZN(n_0_0_222));
   OAI22_X1 i_0_0_296 (.A1(n_0_0_174), .A2(n_0_0_221), .B1(n_0_0_110), .B2(
      n_0_0_222), .ZN(n_0_0_223));
   OAI22_X1 i_0_0_297 (.A1(n_0_0_223), .A2(i[2]), .B1(n_0_0_181), .B2(n_0_0_23), 
      .ZN(n_0_0_224));
   AOI22_X1 i_0_0_298 (.A1(n_0_0_224), .A2(n_0_0_19), .B1(n_0_0_202), .B2(i[1]), 
      .ZN(n_0_0_225));
   OAI22_X1 i_0_0_299 (.A1(n_0_0_213), .A2(n_0_0_15), .B1(n_0_0_225), .B2(i[0]), 
      .ZN(n_0_0_226));
   OAI21_X1 i_0_0_300 (.A(n_0_0_220), .B1(n_0_0_102), .B2(n_0_0_226), .ZN(
      partialProd[13]));
   INV_X1 i_0_0_301 (.A(extended_M[6]), .ZN(n_0_0_227));
   INV_X1 i_0_0_302 (.A(extended_M[14]), .ZN(n_0_0_228));
   OAI22_X1 i_0_0_303 (.A1(n_0_0_174), .A2(n_0_0_227), .B1(n_0_0_110), .B2(
      n_0_0_228), .ZN(n_0_0_229));
   OAI22_X1 i_0_0_304 (.A1(n_0_0_229), .A2(i[2]), .B1(n_0_0_186), .B2(n_0_0_23), 
      .ZN(n_0_0_230));
   AOI22_X1 i_0_0_305 (.A1(n_0_0_207), .A2(i[1]), .B1(n_0_0_230), .B2(n_0_0_19), 
      .ZN(n_0_0_231));
   OAI221_X1 i_0_0_306 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_219), .C1(i[0]), 
      .C2(n_0_0_231), .ZN(n_0_0_232));
   INV_X1 i_0_0_307 (.A(extended_M_mul_neg_one[6]), .ZN(n_0_0_233));
   INV_X1 i_0_0_308 (.A(extended_M_mul_neg_one[14]), .ZN(n_0_0_234));
   OAI22_X1 i_0_0_309 (.A1(n_0_0_174), .A2(n_0_0_233), .B1(n_0_0_110), .B2(
      n_0_0_234), .ZN(n_0_0_235));
   OAI22_X1 i_0_0_310 (.A1(n_0_0_235), .A2(i[2]), .B1(n_0_0_191), .B2(n_0_0_23), 
      .ZN(n_0_0_236));
   AOI22_X1 i_0_0_311 (.A1(n_0_0_212), .A2(i[1]), .B1(n_0_0_236), .B2(n_0_0_19), 
      .ZN(n_0_0_237));
   OAI22_X1 i_0_0_312 (.A1(n_0_0_237), .A2(i[0]), .B1(n_0_0_225), .B2(n_0_0_15), 
      .ZN(n_0_0_238));
   OAI21_X1 i_0_0_313 (.A(n_0_0_232), .B1(n_0_0_102), .B2(n_0_0_238), .ZN(
      partialProd[14]));
   INV_X1 i_0_0_314 (.A(extended_M[7]), .ZN(n_0_0_239));
   INV_X1 i_0_0_315 (.A(extended_M[15]), .ZN(n_0_0_240));
   OAI22_X1 i_0_0_316 (.A1(n_0_0_174), .A2(n_0_0_239), .B1(n_0_0_110), .B2(
      n_0_0_240), .ZN(n_0_0_241));
   OAI22_X1 i_0_0_317 (.A1(n_0_0_241), .A2(i[2]), .B1(n_0_0_196), .B2(n_0_0_23), 
      .ZN(n_0_0_242));
   AOI22_X1 i_0_0_318 (.A1(n_0_0_242), .A2(n_0_0_19), .B1(n_0_0_218), .B2(i[1]), 
      .ZN(n_0_0_243));
   OAI221_X1 i_0_0_319 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_231), .C1(i[0]), 
      .C2(n_0_0_243), .ZN(n_0_0_244));
   INV_X1 i_0_0_320 (.A(extended_M_mul_neg_one[7]), .ZN(n_0_0_245));
   INV_X1 i_0_0_321 (.A(extended_M_mul_neg_one[15]), .ZN(n_0_0_246));
   OAI22_X1 i_0_0_322 (.A1(n_0_0_174), .A2(n_0_0_245), .B1(n_0_0_110), .B2(
      n_0_0_246), .ZN(n_0_0_247));
   OAI22_X1 i_0_0_323 (.A1(n_0_0_247), .A2(i[2]), .B1(n_0_0_201), .B2(n_0_0_23), 
      .ZN(n_0_0_248));
   AOI22_X1 i_0_0_324 (.A1(n_0_0_248), .A2(n_0_0_19), .B1(n_0_0_224), .B2(i[1]), 
      .ZN(n_0_0_249));
   OAI22_X1 i_0_0_325 (.A1(n_0_0_237), .A2(n_0_0_15), .B1(n_0_0_249), .B2(i[0]), 
      .ZN(n_0_0_250));
   OAI21_X1 i_0_0_326 (.A(n_0_0_244), .B1(n_0_0_102), .B2(n_0_0_250), .ZN(
      partialProd[15]));
   NAND2_X1 i_0_0_327 (.A1(extended_M[0]), .A2(i[4]), .ZN(n_0_0_251));
   INV_X1 i_0_0_328 (.A(extended_M[16]), .ZN(n_0_0_252));
   OAI21_X1 i_0_0_329 (.A(n_0_0_251), .B1(n_0_0_252), .B2(i[4]), .ZN(n_0_0_253));
   INV_X1 i_0_0_330 (.A(n_0_0_253), .ZN(n_0_0_254));
   OAI22_X1 i_0_0_331 (.A1(n_0_0_254), .A2(n_0_0_11), .B1(n_0_0_174), .B2(
      n_0_0_164), .ZN(n_0_0_255));
   OAI22_X1 i_0_0_332 (.A1(n_0_0_255), .A2(i[2]), .B1(n_0_0_206), .B2(n_0_0_23), 
      .ZN(n_0_0_256));
   AOI22_X1 i_0_0_333 (.A1(n_0_0_256), .A2(n_0_0_19), .B1(n_0_0_230), .B2(i[1]), 
      .ZN(n_0_0_257));
   OAI221_X1 i_0_0_334 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_243), .C1(i[0]), 
      .C2(n_0_0_257), .ZN(n_0_0_258));
   INV_X1 i_0_0_335 (.A(extended_M_mul_neg_one[16]), .ZN(n_0_0_259));
   OAI21_X1 i_0_0_336 (.A(n_0_0_251), .B1(n_0_0_259), .B2(i[4]), .ZN(n_0_0_260));
   NAND2_X1 i_0_0_337 (.A1(n_0_0_260), .A2(n_0_0_10), .ZN(n_0_0_261));
   OAI22_X1 i_0_0_338 (.A1(n_0_0_261), .A2(i[3]), .B1(n_0_0_174), .B2(n_0_0_169), 
      .ZN(n_0_0_262));
   OAI22_X1 i_0_0_339 (.A1(n_0_0_262), .A2(i[2]), .B1(n_0_0_211), .B2(n_0_0_23), 
      .ZN(n_0_0_263));
   AOI22_X1 i_0_0_340 (.A1(n_0_0_263), .A2(n_0_0_19), .B1(n_0_0_236), .B2(i[1]), 
      .ZN(n_0_0_264));
   OAI22_X1 i_0_0_341 (.A1(n_0_0_264), .A2(i[0]), .B1(n_0_0_249), .B2(n_0_0_15), 
      .ZN(n_0_0_265));
   OAI21_X1 i_0_0_342 (.A(n_0_0_258), .B1(n_0_0_102), .B2(n_0_0_265), .ZN(
      partialProd[16]));
   AOI22_X1 i_0_0_343 (.A1(n_0_0_54), .A2(extended_M[17]), .B1(extended_M[1]), 
      .B2(i[4]), .ZN(n_0_0_266));
   OAI22_X1 i_0_0_344 (.A1(n_0_0_174), .A2(n_0_0_175), .B1(n_0_0_266), .B2(
      n_0_0_11), .ZN(n_0_0_267));
   OAI22_X1 i_0_0_345 (.A1(n_0_0_267), .A2(i[2]), .B1(n_0_0_217), .B2(n_0_0_23), 
      .ZN(n_0_0_268));
   AOI22_X1 i_0_0_346 (.A1(n_0_0_268), .A2(n_0_0_19), .B1(n_0_0_242), .B2(i[1]), 
      .ZN(n_0_0_269));
   OAI221_X1 i_0_0_347 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_257), .C1(i[0]), 
      .C2(n_0_0_269), .ZN(n_0_0_270));
   INV_X1 i_0_0_348 (.A(extended_M_mul_neg_one[17]), .ZN(n_0_0_271));
   AOI22_X1 i_0_0_349 (.A1(n_0_0_271), .A2(n_0_0_54), .B1(n_0_0_108), .B2(i[4]), 
      .ZN(n_0_0_272));
   NAND2_X1 i_0_0_350 (.A1(n_0_0_272), .A2(n_0_0_10), .ZN(n_0_0_273));
   OAI22_X1 i_0_0_351 (.A1(n_0_0_273), .A2(i[3]), .B1(n_0_0_174), .B2(n_0_0_180), 
      .ZN(n_0_0_274));
   OAI22_X1 i_0_0_352 (.A1(n_0_0_274), .A2(i[2]), .B1(n_0_0_223), .B2(n_0_0_23), 
      .ZN(n_0_0_275));
   AOI22_X1 i_0_0_353 (.A1(n_0_0_275), .A2(n_0_0_19), .B1(n_0_0_248), .B2(i[1]), 
      .ZN(n_0_0_276));
   OAI22_X1 i_0_0_354 (.A1(n_0_0_264), .A2(n_0_0_15), .B1(n_0_0_276), .B2(i[0]), 
      .ZN(n_0_0_277));
   OAI21_X1 i_0_0_355 (.A(n_0_0_270), .B1(n_0_0_102), .B2(n_0_0_277), .ZN(
      partialProd[17]));
   AOI22_X1 i_0_0_356 (.A1(n_0_0_54), .A2(extended_M[18]), .B1(extended_M[2]), 
      .B2(i[4]), .ZN(n_0_0_278));
   OAI22_X1 i_0_0_357 (.A1(n_0_0_174), .A2(n_0_0_185), .B1(n_0_0_278), .B2(
      n_0_0_11), .ZN(n_0_0_279));
   OAI22_X1 i_0_0_358 (.A1(n_0_0_279), .A2(i[2]), .B1(n_0_0_229), .B2(n_0_0_23), 
      .ZN(n_0_0_280));
   AOI22_X1 i_0_0_359 (.A1(n_0_0_256), .A2(i[1]), .B1(n_0_0_280), .B2(n_0_0_19), 
      .ZN(n_0_0_281));
   OAI221_X1 i_0_0_360 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_269), .C1(i[0]), 
      .C2(n_0_0_281), .ZN(n_0_0_282));
   AOI22_X1 i_0_0_361 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[18]), .B1(
      extended_M_mul_neg_one[2]), .B2(i[4]), .ZN(n_0_0_283));
   OAI22_X1 i_0_0_362 (.A1(n_0_0_174), .A2(n_0_0_190), .B1(n_0_0_283), .B2(
      n_0_0_11), .ZN(n_0_0_284));
   OAI22_X1 i_0_0_363 (.A1(n_0_0_284), .A2(i[2]), .B1(n_0_0_235), .B2(n_0_0_23), 
      .ZN(n_0_0_285));
   AOI22_X1 i_0_0_364 (.A1(n_0_0_263), .A2(i[1]), .B1(n_0_0_285), .B2(n_0_0_19), 
      .ZN(n_0_0_286));
   OAI22_X1 i_0_0_365 (.A1(n_0_0_286), .A2(i[0]), .B1(n_0_0_276), .B2(n_0_0_15), 
      .ZN(n_0_0_287));
   OAI21_X1 i_0_0_366 (.A(n_0_0_282), .B1(n_0_0_102), .B2(n_0_0_287), .ZN(
      partialProd[18]));
   AOI22_X1 i_0_0_367 (.A1(n_0_0_54), .A2(extended_M[19]), .B1(extended_M[3]), 
      .B2(i[4]), .ZN(n_0_0_288));
   OAI22_X1 i_0_0_368 (.A1(n_0_0_174), .A2(n_0_0_195), .B1(n_0_0_288), .B2(
      n_0_0_11), .ZN(n_0_0_289));
   OAI22_X1 i_0_0_369 (.A1(n_0_0_289), .A2(i[2]), .B1(n_0_0_241), .B2(n_0_0_23), 
      .ZN(n_0_0_290));
   AOI22_X1 i_0_0_370 (.A1(n_0_0_290), .A2(n_0_0_19), .B1(n_0_0_268), .B2(i[1]), 
      .ZN(n_0_0_291));
   OAI221_X1 i_0_0_371 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_281), .C1(i[0]), 
      .C2(n_0_0_291), .ZN(n_0_0_292));
   AOI22_X1 i_0_0_372 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[19]), .B1(
      extended_M_mul_neg_one[3]), .B2(i[4]), .ZN(n_0_0_293));
   OAI22_X1 i_0_0_373 (.A1(n_0_0_174), .A2(n_0_0_200), .B1(n_0_0_293), .B2(
      n_0_0_11), .ZN(n_0_0_294));
   OAI22_X1 i_0_0_374 (.A1(n_0_0_294), .A2(i[2]), .B1(n_0_0_247), .B2(n_0_0_23), 
      .ZN(n_0_0_295));
   AOI22_X1 i_0_0_375 (.A1(n_0_0_275), .A2(i[1]), .B1(n_0_0_295), .B2(n_0_0_19), 
      .ZN(n_0_0_296));
   OAI22_X1 i_0_0_376 (.A1(n_0_0_286), .A2(n_0_0_15), .B1(n_0_0_296), .B2(i[0]), 
      .ZN(n_0_0_297));
   OAI21_X1 i_0_0_377 (.A(n_0_0_292), .B1(n_0_0_102), .B2(n_0_0_297), .ZN(
      partialProd[19]));
   AOI22_X1 i_0_0_378 (.A1(n_0_0_54), .A2(extended_M[20]), .B1(extended_M[4]), 
      .B2(i[4]), .ZN(n_0_0_298));
   OAI22_X1 i_0_0_379 (.A1(n_0_0_174), .A2(n_0_0_205), .B1(n_0_0_298), .B2(
      n_0_0_11), .ZN(n_0_0_299));
   OAI22_X1 i_0_0_380 (.A1(n_0_0_255), .A2(n_0_0_23), .B1(n_0_0_299), .B2(i[2]), 
      .ZN(n_0_0_300));
   AOI22_X1 i_0_0_381 (.A1(n_0_0_300), .A2(n_0_0_19), .B1(n_0_0_280), .B2(i[1]), 
      .ZN(n_0_0_301));
   OAI221_X1 i_0_0_382 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_291), .C1(i[0]), 
      .C2(n_0_0_301), .ZN(n_0_0_302));
   AOI22_X1 i_0_0_383 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[20]), .B1(
      extended_M_mul_neg_one[4]), .B2(i[4]), .ZN(n_0_0_303));
   OAI22_X1 i_0_0_384 (.A1(n_0_0_174), .A2(n_0_0_210), .B1(n_0_0_303), .B2(
      n_0_0_11), .ZN(n_0_0_304));
   OAI22_X1 i_0_0_385 (.A1(n_0_0_262), .A2(n_0_0_23), .B1(n_0_0_304), .B2(i[2]), 
      .ZN(n_0_0_305));
   AOI22_X1 i_0_0_386 (.A1(n_0_0_305), .A2(n_0_0_19), .B1(n_0_0_285), .B2(i[1]), 
      .ZN(n_0_0_306));
   OAI22_X1 i_0_0_387 (.A1(n_0_0_306), .A2(i[0]), .B1(n_0_0_296), .B2(n_0_0_15), 
      .ZN(n_0_0_307));
   OAI21_X1 i_0_0_388 (.A(n_0_0_302), .B1(n_0_0_102), .B2(n_0_0_307), .ZN(
      partialProd[20]));
   AOI22_X1 i_0_0_389 (.A1(n_0_0_54), .A2(extended_M[21]), .B1(extended_M[5]), 
      .B2(i[4]), .ZN(n_0_0_308));
   OAI22_X1 i_0_0_390 (.A1(n_0_0_174), .A2(n_0_0_216), .B1(n_0_0_308), .B2(
      n_0_0_11), .ZN(n_0_0_309));
   OAI22_X1 i_0_0_391 (.A1(n_0_0_267), .A2(n_0_0_23), .B1(n_0_0_309), .B2(i[2]), 
      .ZN(n_0_0_310));
   AOI22_X1 i_0_0_392 (.A1(n_0_0_290), .A2(i[1]), .B1(n_0_0_310), .B2(n_0_0_19), 
      .ZN(n_0_0_311));
   OAI221_X1 i_0_0_393 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_301), .C1(i[0]), 
      .C2(n_0_0_311), .ZN(n_0_0_312));
   AOI22_X1 i_0_0_394 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[21]), .B1(
      extended_M_mul_neg_one[5]), .B2(i[4]), .ZN(n_0_0_313));
   OAI22_X1 i_0_0_395 (.A1(n_0_0_174), .A2(n_0_0_222), .B1(n_0_0_313), .B2(
      n_0_0_11), .ZN(n_0_0_314));
   OAI22_X1 i_0_0_396 (.A1(n_0_0_314), .A2(i[2]), .B1(n_0_0_274), .B2(n_0_0_23), 
      .ZN(n_0_0_315));
   AOI22_X1 i_0_0_397 (.A1(n_0_0_315), .A2(n_0_0_19), .B1(n_0_0_295), .B2(i[1]), 
      .ZN(n_0_0_316));
   OAI22_X1 i_0_0_398 (.A1(n_0_0_306), .A2(n_0_0_15), .B1(n_0_0_316), .B2(i[0]), 
      .ZN(n_0_0_317));
   OAI21_X1 i_0_0_399 (.A(n_0_0_312), .B1(n_0_0_102), .B2(n_0_0_317), .ZN(
      partialProd[21]));
   AOI22_X1 i_0_0_400 (.A1(n_0_0_54), .A2(extended_M[22]), .B1(extended_M[6]), 
      .B2(i[4]), .ZN(n_0_0_318));
   OAI22_X1 i_0_0_401 (.A1(n_0_0_174), .A2(n_0_0_228), .B1(n_0_0_318), .B2(
      n_0_0_11), .ZN(n_0_0_319));
   OAI22_X1 i_0_0_402 (.A1(n_0_0_319), .A2(i[2]), .B1(n_0_0_279), .B2(n_0_0_23), 
      .ZN(n_0_0_320));
   AOI22_X1 i_0_0_403 (.A1(n_0_0_300), .A2(i[1]), .B1(n_0_0_320), .B2(n_0_0_19), 
      .ZN(n_0_0_321));
   OAI221_X1 i_0_0_404 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_311), .C1(i[0]), 
      .C2(n_0_0_321), .ZN(n_0_0_322));
   AOI22_X1 i_0_0_405 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[22]), .B1(
      extended_M_mul_neg_one[6]), .B2(i[4]), .ZN(n_0_0_323));
   OAI22_X1 i_0_0_406 (.A1(n_0_0_174), .A2(n_0_0_234), .B1(n_0_0_323), .B2(
      n_0_0_11), .ZN(n_0_0_324));
   OAI22_X1 i_0_0_407 (.A1(n_0_0_284), .A2(n_0_0_23), .B1(n_0_0_324), .B2(i[2]), 
      .ZN(n_0_0_325));
   AOI22_X1 i_0_0_408 (.A1(n_0_0_305), .A2(i[1]), .B1(n_0_0_325), .B2(n_0_0_19), 
      .ZN(n_0_0_326));
   OAI22_X1 i_0_0_409 (.A1(n_0_0_326), .A2(i[0]), .B1(n_0_0_316), .B2(n_0_0_15), 
      .ZN(n_0_0_327));
   OAI21_X1 i_0_0_410 (.A(n_0_0_322), .B1(n_0_0_102), .B2(n_0_0_327), .ZN(
      partialProd[22]));
   AOI22_X1 i_0_0_411 (.A1(n_0_0_54), .A2(extended_M[23]), .B1(extended_M[7]), 
      .B2(i[4]), .ZN(n_0_0_328));
   OAI22_X1 i_0_0_412 (.A1(n_0_0_174), .A2(n_0_0_240), .B1(n_0_0_328), .B2(
      n_0_0_11), .ZN(n_0_0_329));
   OAI22_X1 i_0_0_413 (.A1(n_0_0_289), .A2(n_0_0_23), .B1(n_0_0_329), .B2(i[2]), 
      .ZN(n_0_0_330));
   AOI22_X1 i_0_0_414 (.A1(n_0_0_330), .A2(n_0_0_19), .B1(n_0_0_310), .B2(i[1]), 
      .ZN(n_0_0_331));
   OAI221_X1 i_0_0_415 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_321), .C1(i[0]), 
      .C2(n_0_0_331), .ZN(n_0_0_332));
   AOI22_X1 i_0_0_416 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[23]), .B1(
      extended_M_mul_neg_one[7]), .B2(i[4]), .ZN(n_0_0_333));
   OAI22_X1 i_0_0_417 (.A1(n_0_0_174), .A2(n_0_0_246), .B1(n_0_0_333), .B2(
      n_0_0_11), .ZN(n_0_0_334));
   OAI22_X1 i_0_0_418 (.A1(n_0_0_294), .A2(n_0_0_23), .B1(n_0_0_334), .B2(i[2]), 
      .ZN(n_0_0_335));
   AOI22_X1 i_0_0_419 (.A1(n_0_0_315), .A2(i[1]), .B1(n_0_0_335), .B2(n_0_0_19), 
      .ZN(n_0_0_336));
   OAI22_X1 i_0_0_420 (.A1(n_0_0_336), .A2(i[0]), .B1(n_0_0_326), .B2(n_0_0_15), 
      .ZN(n_0_0_337));
   OAI21_X1 i_0_0_421 (.A(n_0_0_332), .B1(n_0_0_102), .B2(n_0_0_337), .ZN(
      partialProd[23]));
   OAI22_X1 i_0_0_422 (.A1(n_0_0_54), .A2(extended_M[8]), .B1(extended_M[24]), 
      .B2(i[4]), .ZN(n_0_0_338));
   INV_X1 i_0_0_423 (.A(n_0_0_338), .ZN(n_0_0_339));
   AOI22_X1 i_0_0_424 (.A1(n_0_0_253), .A2(i[3]), .B1(n_0_0_339), .B2(n_0_0_9), 
      .ZN(n_0_0_340));
   NOR2_X1 i_0_0_425 (.A1(n_0_0_340), .A2(i[5]), .ZN(n_0_0_341));
   OAI22_X1 i_0_0_426 (.A1(n_0_0_341), .A2(i[2]), .B1(n_0_0_299), .B2(n_0_0_23), 
      .ZN(n_0_0_342));
   AOI22_X1 i_0_0_427 (.A1(n_0_0_342), .A2(n_0_0_19), .B1(n_0_0_320), .B2(i[1]), 
      .ZN(n_0_0_343));
   OAI221_X1 i_0_0_428 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_331), .C1(i[0]), 
      .C2(n_0_0_343), .ZN(n_0_0_344));
   OAI22_X1 i_0_0_429 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[8]), .B1(
      extended_M_mul_neg_one[24]), .B2(i[4]), .ZN(n_0_0_345));
   OAI22_X1 i_0_0_430 (.A1(n_0_0_261), .A2(n_0_0_9), .B1(n_0_0_345), .B2(
      n_0_0_11), .ZN(n_0_0_346));
   OAI22_X1 i_0_0_431 (.A1(n_0_0_346), .A2(i[2]), .B1(n_0_0_304), .B2(n_0_0_23), 
      .ZN(n_0_0_347));
   AOI22_X1 i_0_0_432 (.A1(n_0_0_347), .A2(n_0_0_19), .B1(n_0_0_325), .B2(i[1]), 
      .ZN(n_0_0_348));
   OAI22_X1 i_0_0_433 (.A1(n_0_0_336), .A2(n_0_0_15), .B1(n_0_0_348), .B2(i[0]), 
      .ZN(n_0_0_349));
   OAI21_X1 i_0_0_434 (.A(n_0_0_344), .B1(n_0_0_102), .B2(n_0_0_349), .ZN(
      partialProd[24]));
   AOI22_X1 i_0_0_435 (.A1(n_0_0_54), .A2(extended_M[25]), .B1(extended_M[9]), 
      .B2(i[4]), .ZN(n_0_0_350));
   OAI22_X1 i_0_0_436 (.A1(n_0_0_350), .A2(n_0_0_11), .B1(n_0_0_266), .B2(
      n_0_0_161), .ZN(n_0_0_351));
   OAI22_X1 i_0_0_437 (.A1(n_0_0_309), .A2(n_0_0_23), .B1(n_0_0_351), .B2(i[2]), 
      .ZN(n_0_0_352));
   AOI22_X1 i_0_0_438 (.A1(n_0_0_330), .A2(i[1]), .B1(n_0_0_352), .B2(n_0_0_19), 
      .ZN(n_0_0_353));
   OAI221_X1 i_0_0_439 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_343), .C1(i[0]), 
      .C2(n_0_0_353), .ZN(n_0_0_354));
   AOI22_X1 i_0_0_440 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[25]), .B1(
      extended_M_mul_neg_one[9]), .B2(i[4]), .ZN(n_0_0_355));
   OAI22_X1 i_0_0_441 (.A1(n_0_0_273), .A2(n_0_0_9), .B1(n_0_0_355), .B2(
      n_0_0_11), .ZN(n_0_0_356));
   OAI22_X1 i_0_0_442 (.A1(n_0_0_356), .A2(i[2]), .B1(n_0_0_314), .B2(n_0_0_23), 
      .ZN(n_0_0_357));
   AOI22_X1 i_0_0_443 (.A1(n_0_0_357), .A2(n_0_0_19), .B1(n_0_0_335), .B2(i[1]), 
      .ZN(n_0_0_358));
   OAI22_X1 i_0_0_444 (.A1(n_0_0_358), .A2(i[0]), .B1(n_0_0_348), .B2(n_0_0_15), 
      .ZN(n_0_0_359));
   OAI21_X1 i_0_0_445 (.A(n_0_0_354), .B1(n_0_0_102), .B2(n_0_0_359), .ZN(
      partialProd[25]));
   AOI22_X1 i_0_0_446 (.A1(n_0_0_54), .A2(extended_M[26]), .B1(extended_M[10]), 
      .B2(i[4]), .ZN(n_0_0_360));
   OAI22_X1 i_0_0_447 (.A1(n_0_0_360), .A2(n_0_0_11), .B1(n_0_0_278), .B2(
      n_0_0_161), .ZN(n_0_0_361));
   OAI22_X1 i_0_0_448 (.A1(n_0_0_319), .A2(n_0_0_23), .B1(n_0_0_361), .B2(i[2]), 
      .ZN(n_0_0_362));
   AOI22_X1 i_0_0_449 (.A1(n_0_0_342), .A2(i[1]), .B1(n_0_0_362), .B2(n_0_0_19), 
      .ZN(n_0_0_363));
   OAI221_X1 i_0_0_450 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_353), .C1(i[0]), 
      .C2(n_0_0_363), .ZN(n_0_0_364));
   OAI22_X1 i_0_0_451 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[10]), .B1(
      extended_M_mul_neg_one[26]), .B2(i[4]), .ZN(n_0_0_365));
   OR2_X1 i_0_0_452 (.A1(n_0_0_365), .A2(i[5]), .ZN(n_0_0_366));
   OAI22_X1 i_0_0_453 (.A1(n_0_0_366), .A2(i[3]), .B1(n_0_0_283), .B2(n_0_0_161), 
      .ZN(n_0_0_367));
   OAI22_X1 i_0_0_454 (.A1(n_0_0_367), .A2(i[2]), .B1(n_0_0_324), .B2(n_0_0_23), 
      .ZN(n_0_0_368));
   AOI22_X1 i_0_0_455 (.A1(n_0_0_368), .A2(n_0_0_19), .B1(n_0_0_347), .B2(i[1]), 
      .ZN(n_0_0_369));
   OAI22_X1 i_0_0_456 (.A1(n_0_0_358), .A2(n_0_0_15), .B1(n_0_0_369), .B2(i[0]), 
      .ZN(n_0_0_370));
   OAI21_X1 i_0_0_457 (.A(n_0_0_364), .B1(n_0_0_102), .B2(n_0_0_370), .ZN(
      partialProd[26]));
   AOI22_X1 i_0_0_458 (.A1(n_0_0_54), .A2(extended_M[27]), .B1(extended_M[11]), 
      .B2(i[4]), .ZN(n_0_0_371));
   OAI22_X1 i_0_0_459 (.A1(n_0_0_371), .A2(n_0_0_11), .B1(n_0_0_288), .B2(
      n_0_0_161), .ZN(n_0_0_372));
   OAI22_X1 i_0_0_460 (.A1(n_0_0_329), .A2(n_0_0_23), .B1(n_0_0_372), .B2(i[2]), 
      .ZN(n_0_0_373));
   AOI22_X1 i_0_0_461 (.A1(n_0_0_373), .A2(n_0_0_19), .B1(n_0_0_352), .B2(i[1]), 
      .ZN(n_0_0_374));
   OAI221_X1 i_0_0_462 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_363), .C1(i[0]), 
      .C2(n_0_0_374), .ZN(n_0_0_375));
   INV_X1 i_0_0_463 (.A(extended_M_mul_neg_one[27]), .ZN(n_0_0_376));
   AOI22_X1 i_0_0_464 (.A1(n_0_0_376), .A2(n_0_0_54), .B1(n_0_0_200), .B2(i[4]), 
      .ZN(n_0_0_377));
   NAND2_X1 i_0_0_465 (.A1(n_0_0_377), .A2(n_0_0_10), .ZN(n_0_0_378));
   OAI22_X1 i_0_0_466 (.A1(n_0_0_378), .A2(i[3]), .B1(n_0_0_293), .B2(n_0_0_161), 
      .ZN(n_0_0_379));
   OAI22_X1 i_0_0_467 (.A1(n_0_0_379), .A2(i[2]), .B1(n_0_0_334), .B2(n_0_0_23), 
      .ZN(n_0_0_380));
   AOI22_X1 i_0_0_468 (.A1(n_0_0_357), .A2(i[1]), .B1(n_0_0_380), .B2(n_0_0_19), 
      .ZN(n_0_0_381));
   OAI22_X1 i_0_0_469 (.A1(n_0_0_381), .A2(i[0]), .B1(n_0_0_369), .B2(n_0_0_15), 
      .ZN(n_0_0_382));
   OAI21_X1 i_0_0_470 (.A(n_0_0_375), .B1(n_0_0_102), .B2(n_0_0_382), .ZN(
      partialProd[27]));
   AOI22_X1 i_0_0_471 (.A1(n_0_0_54), .A2(extended_M[28]), .B1(extended_M[12]), 
      .B2(i[4]), .ZN(n_0_0_383));
   INV_X1 i_0_0_472 (.A(n_0_0_383), .ZN(n_0_0_384));
   INV_X1 i_0_0_473 (.A(n_0_0_298), .ZN(n_0_0_385));
   OAI22_X1 i_0_0_474 (.A1(n_0_0_384), .A2(i[3]), .B1(n_0_0_385), .B2(n_0_0_9), 
      .ZN(n_0_0_386));
   NOR2_X1 i_0_0_475 (.A1(n_0_0_386), .A2(i[5]), .ZN(n_0_0_387));
   OAI22_X1 i_0_0_476 (.A1(n_0_0_341), .A2(n_0_0_23), .B1(n_0_0_387), .B2(i[2]), 
      .ZN(n_0_0_388));
   AOI22_X1 i_0_0_477 (.A1(n_0_0_388), .A2(n_0_0_19), .B1(i[1]), .B2(n_0_0_362), 
      .ZN(n_0_0_389));
   OAI221_X1 i_0_0_478 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_374), .C1(i[0]), 
      .C2(n_0_0_389), .ZN(n_0_0_390));
   AOI22_X1 i_0_0_479 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[28]), .B1(
      extended_M_mul_neg_one[12]), .B2(i[4]), .ZN(n_0_0_391));
   OAI22_X1 i_0_0_480 (.A1(n_0_0_391), .A2(i[3]), .B1(n_0_0_303), .B2(n_0_0_9), 
      .ZN(n_0_0_392));
   AND2_X1 i_0_0_481 (.A1(n_0_0_392), .A2(n_0_0_10), .ZN(n_0_0_393));
   OAI22_X1 i_0_0_482 (.A1(n_0_0_393), .A2(i[2]), .B1(n_0_0_346), .B2(n_0_0_23), 
      .ZN(n_0_0_394));
   AOI22_X1 i_0_0_483 (.A1(n_0_0_394), .A2(n_0_0_19), .B1(n_0_0_368), .B2(i[1]), 
      .ZN(n_0_0_395));
   OAI22_X1 i_0_0_484 (.A1(n_0_0_381), .A2(n_0_0_15), .B1(n_0_0_395), .B2(i[0]), 
      .ZN(n_0_0_396));
   OAI21_X1 i_0_0_485 (.A(n_0_0_390), .B1(n_0_0_102), .B2(n_0_0_396), .ZN(
      partialProd[28]));
   AOI22_X1 i_0_0_486 (.A1(n_0_0_54), .A2(extended_M[29]), .B1(extended_M[13]), 
      .B2(i[4]), .ZN(n_0_0_397));
   OAI22_X1 i_0_0_487 (.A1(n_0_0_397), .A2(n_0_0_11), .B1(n_0_0_308), .B2(
      n_0_0_161), .ZN(n_0_0_398));
   OAI22_X1 i_0_0_488 (.A1(n_0_0_351), .A2(n_0_0_23), .B1(n_0_0_398), .B2(i[2]), 
      .ZN(n_0_0_399));
   AOI22_X1 i_0_0_489 (.A1(n_0_0_373), .A2(i[1]), .B1(n_0_0_399), .B2(n_0_0_19), 
      .ZN(n_0_0_400));
   OAI221_X1 i_0_0_490 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_389), .C1(i[0]), 
      .C2(n_0_0_400), .ZN(n_0_0_401));
   AOI22_X1 i_0_0_491 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[29]), .B1(
      extended_M_mul_neg_one[13]), .B2(i[4]), .ZN(n_0_0_402));
   INV_X1 i_0_0_492 (.A(n_0_0_402), .ZN(n_0_0_403));
   INV_X1 i_0_0_493 (.A(n_0_0_313), .ZN(n_0_0_404));
   AOI22_X1 i_0_0_494 (.A1(n_0_0_403), .A2(n_0_0_9), .B1(n_0_0_404), .B2(i[3]), 
      .ZN(n_0_0_405));
   NOR2_X1 i_0_0_495 (.A1(n_0_0_405), .A2(i[5]), .ZN(n_0_0_406));
   OAI22_X1 i_0_0_496 (.A1(n_0_0_406), .A2(i[2]), .B1(n_0_0_356), .B2(n_0_0_23), 
      .ZN(n_0_0_407));
   AOI22_X1 i_0_0_497 (.A1(n_0_0_407), .A2(n_0_0_19), .B1(n_0_0_380), .B2(i[1]), 
      .ZN(n_0_0_408));
   OAI22_X1 i_0_0_498 (.A1(n_0_0_395), .A2(n_0_0_15), .B1(n_0_0_408), .B2(i[0]), 
      .ZN(n_0_0_409));
   OAI21_X1 i_0_0_499 (.A(n_0_0_401), .B1(n_0_0_102), .B2(n_0_0_409), .ZN(
      partialProd[29]));
   INV_X1 i_0_0_500 (.A(n_0_0_318), .ZN(n_0_0_410));
   AOI22_X1 i_0_0_501 (.A1(n_0_0_54), .A2(extended_M[30]), .B1(extended_M[14]), 
      .B2(i[4]), .ZN(n_0_0_411));
   INV_X1 i_0_0_502 (.A(n_0_0_411), .ZN(n_0_0_412));
   OAI22_X1 i_0_0_503 (.A1(n_0_0_410), .A2(n_0_0_9), .B1(n_0_0_412), .B2(i[3]), 
      .ZN(n_0_0_413));
   NOR2_X1 i_0_0_504 (.A1(n_0_0_413), .A2(i[5]), .ZN(n_0_0_414));
   OAI22_X1 i_0_0_505 (.A1(n_0_0_414), .A2(i[2]), .B1(n_0_0_361), .B2(n_0_0_23), 
      .ZN(n_0_0_415));
   AOI22_X1 i_0_0_506 (.A1(n_0_0_388), .A2(i[1]), .B1(n_0_0_415), .B2(n_0_0_19), 
      .ZN(n_0_0_416));
   OAI221_X1 i_0_0_507 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_400), .C1(i[0]), 
      .C2(n_0_0_416), .ZN(n_0_0_417));
   OAI22_X1 i_0_0_508 (.A1(n_0_0_54), .A2(extended_M_mul_neg_one[14]), .B1(
      extended_M_mul_neg_one[30]), .B2(i[4]), .ZN(n_0_0_418));
   OAI22_X1 i_0_0_509 (.A1(n_0_0_418), .A2(i[3]), .B1(n_0_0_323), .B2(n_0_0_9), 
      .ZN(n_0_0_419));
   AND2_X1 i_0_0_510 (.A1(n_0_0_419), .A2(n_0_0_10), .ZN(n_0_0_420));
   OAI22_X1 i_0_0_511 (.A1(n_0_0_420), .A2(i[2]), .B1(n_0_0_367), .B2(n_0_0_23), 
      .ZN(n_0_0_421));
   AOI22_X1 i_0_0_512 (.A1(n_0_0_421), .A2(n_0_0_19), .B1(n_0_0_394), .B2(i[1]), 
      .ZN(n_0_0_422));
   OAI22_X1 i_0_0_513 (.A1(n_0_0_422), .A2(i[0]), .B1(n_0_0_408), .B2(n_0_0_15), 
      .ZN(n_0_0_423));
   OAI21_X1 i_0_0_514 (.A(n_0_0_417), .B1(n_0_0_102), .B2(n_0_0_423), .ZN(
      partialProd[30]));
   NAND2_X1 i_0_0_515 (.A1(n_0_0_10), .A2(extended_M[63]), .ZN(n_0_0_424));
   NOR2_X1 i_0_0_516 (.A1(n_0_0_424), .A2(i[4]), .ZN(n_0_0_425));
   NOR2_X1 i_0_0_517 (.A1(n_0_0_54), .A2(i[5]), .ZN(n_0_0_426));
   AOI21_X1 i_0_0_518 (.A(n_0_0_425), .B1(extended_M[15]), .B2(n_0_0_426), 
      .ZN(n_0_0_427));
   OAI22_X1 i_0_0_519 (.A1(n_0_0_427), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_328), 
      .ZN(n_0_0_428));
   OAI22_X1 i_0_0_520 (.A1(n_0_0_428), .A2(i[2]), .B1(n_0_0_23), .B2(n_0_0_372), 
      .ZN(n_0_0_429));
   AOI22_X1 i_0_0_521 (.A1(n_0_0_429), .A2(n_0_0_19), .B1(i[1]), .B2(n_0_0_399), 
      .ZN(n_0_0_430));
   OAI221_X1 i_0_0_522 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_416), .C1(i[0]), 
      .C2(n_0_0_430), .ZN(n_0_0_431));
   NAND2_X1 i_0_0_523 (.A1(n_0_0_10), .A2(extended_M_mul_neg_one[63]), .ZN(
      n_0_0_432));
   NOR2_X1 i_0_0_524 (.A1(n_0_0_432), .A2(i[4]), .ZN(n_0_0_433));
   AOI21_X1 i_0_0_525 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[15]), .B2(
      n_0_0_426), .ZN(n_0_0_434));
   OAI22_X1 i_0_0_526 (.A1(n_0_0_434), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_333), 
      .ZN(n_0_0_435));
   OAI22_X1 i_0_0_527 (.A1(n_0_0_435), .A2(i[2]), .B1(n_0_0_379), .B2(n_0_0_23), 
      .ZN(n_0_0_436));
   AOI22_X1 i_0_0_528 (.A1(n_0_0_436), .A2(n_0_0_19), .B1(n_0_0_407), .B2(i[1]), 
      .ZN(n_0_0_437));
   OAI22_X1 i_0_0_529 (.A1(n_0_0_437), .A2(i[0]), .B1(n_0_0_422), .B2(n_0_0_15), 
      .ZN(n_0_0_438));
   OAI21_X1 i_0_0_530 (.A(n_0_0_431), .B1(n_0_0_102), .B2(n_0_0_438), .ZN(
      partialProd[31]));
   NOR2_X1 i_0_0_531 (.A1(n_0_0_10), .A2(i[4]), .ZN(n_0_0_439));
   AND2_X1 i_0_0_532 (.A1(n_0_0_439), .A2(extended_M[0]), .ZN(n_0_0_440));
   AOI211_X1 i_0_0_533 (.A(n_0_0_425), .B(n_0_0_440), .C1(extended_M[16]), 
      .C2(n_0_0_426), .ZN(n_0_0_441));
   OAI22_X1 i_0_0_534 (.A1(n_0_0_441), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_338), 
      .ZN(n_0_0_442));
   AOI22_X1 i_0_0_535 (.A1(n_0_0_442), .A2(n_0_0_23), .B1(i[2]), .B2(n_0_0_387), 
      .ZN(n_0_0_443));
   OAI22_X1 i_0_0_536 (.A1(n_0_0_443), .A2(i[1]), .B1(n_0_0_19), .B2(n_0_0_415), 
      .ZN(n_0_0_444));
   OAI221_X1 i_0_0_537 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_430), .C1(i[0]), 
      .C2(n_0_0_444), .ZN(n_0_0_445));
   AOI211_X1 i_0_0_538 (.A(n_0_0_433), .B(n_0_0_440), .C1(
      extended_M_mul_neg_one[16]), .C2(n_0_0_426), .ZN(n_0_0_446));
   OAI22_X1 i_0_0_539 (.A1(n_0_0_446), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_345), 
      .ZN(n_0_0_447));
   AOI22_X1 i_0_0_540 (.A1(n_0_0_447), .A2(n_0_0_23), .B1(i[2]), .B2(n_0_0_393), 
      .ZN(n_0_0_448));
   OAI22_X1 i_0_0_541 (.A1(n_0_0_448), .A2(i[1]), .B1(n_0_0_19), .B2(n_0_0_421), 
      .ZN(n_0_0_449));
   OAI22_X1 i_0_0_542 (.A1(n_0_0_449), .A2(i[0]), .B1(n_0_0_437), .B2(n_0_0_15), 
      .ZN(n_0_0_450));
   OAI21_X1 i_0_0_543 (.A(n_0_0_445), .B1(n_0_0_102), .B2(n_0_0_450), .ZN(
      partialProd[32]));
   AOI221_X1 i_0_0_544 (.A(n_0_0_425), .B1(extended_M[1]), .B2(n_0_0_439), 
      .C1(extended_M[17]), .C2(n_0_0_426), .ZN(n_0_0_451));
   OAI22_X1 i_0_0_545 (.A1(n_0_0_451), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_350), 
      .ZN(n_0_0_452));
   OAI22_X1 i_0_0_546 (.A1(n_0_0_452), .A2(i[2]), .B1(n_0_0_23), .B2(n_0_0_398), 
      .ZN(n_0_0_453));
   AOI22_X1 i_0_0_547 (.A1(n_0_0_453), .A2(n_0_0_19), .B1(n_0_0_429), .B2(i[1]), 
      .ZN(n_0_0_454));
   OAI221_X1 i_0_0_548 (.A(n_0_0_100), .B1(i[0]), .B2(n_0_0_454), .C1(n_0_0_15), 
      .C2(n_0_0_444), .ZN(n_0_0_455));
   AOI221_X1 i_0_0_549 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[17]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[1]), .C2(n_0_0_439), .ZN(n_0_0_456));
   OAI22_X1 i_0_0_550 (.A1(n_0_0_456), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_355), 
      .ZN(n_0_0_457));
   OAI22_X1 i_0_0_551 (.A1(n_0_0_457), .A2(i[2]), .B1(n_0_0_23), .B2(n_0_0_406), 
      .ZN(n_0_0_458));
   AOI22_X1 i_0_0_552 (.A1(n_0_0_458), .A2(n_0_0_19), .B1(i[1]), .B2(n_0_0_436), 
      .ZN(n_0_0_459));
   OAI22_X1 i_0_0_553 (.A1(n_0_0_449), .A2(n_0_0_15), .B1(n_0_0_459), .B2(i[0]), 
      .ZN(n_0_0_460));
   OAI21_X1 i_0_0_554 (.A(n_0_0_455), .B1(n_0_0_102), .B2(n_0_0_460), .ZN(
      partialProd[33]));
   AOI221_X1 i_0_0_555 (.A(n_0_0_425), .B1(extended_M[2]), .B2(n_0_0_439), 
      .C1(extended_M[18]), .C2(n_0_0_426), .ZN(n_0_0_461));
   OAI22_X1 i_0_0_556 (.A1(n_0_0_461), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_360), 
      .ZN(n_0_0_462));
   OAI22_X1 i_0_0_557 (.A1(n_0_0_462), .A2(i[2]), .B1(n_0_0_23), .B2(n_0_0_414), 
      .ZN(n_0_0_463));
   OAI22_X1 i_0_0_558 (.A1(n_0_0_463), .A2(i[1]), .B1(n_0_0_443), .B2(n_0_0_19), 
      .ZN(n_0_0_464));
   OAI221_X1 i_0_0_559 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_454), .C1(i[0]), 
      .C2(n_0_0_464), .ZN(n_0_0_465));
   AOI221_X1 i_0_0_560 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[18]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[2]), .C2(n_0_0_439), .ZN(n_0_0_466));
   OAI22_X1 i_0_0_561 (.A1(n_0_0_466), .A2(i[3]), .B1(n_0_0_9), .B2(n_0_0_366), 
      .ZN(n_0_0_467));
   OAI22_X1 i_0_0_562 (.A1(n_0_0_467), .A2(i[2]), .B1(n_0_0_23), .B2(n_0_0_420), 
      .ZN(n_0_0_468));
   OAI22_X1 i_0_0_563 (.A1(n_0_0_468), .A2(i[1]), .B1(n_0_0_448), .B2(n_0_0_19), 
      .ZN(n_0_0_469));
   OAI22_X1 i_0_0_564 (.A1(n_0_0_469), .A2(i[0]), .B1(n_0_0_459), .B2(n_0_0_15), 
      .ZN(n_0_0_470));
   OAI21_X1 i_0_0_565 (.A(n_0_0_465), .B1(n_0_0_102), .B2(n_0_0_470), .ZN(
      partialProd[34]));
   AOI221_X1 i_0_0_566 (.A(n_0_0_425), .B1(extended_M[3]), .B2(n_0_0_439), 
      .C1(extended_M[19]), .C2(n_0_0_426), .ZN(n_0_0_471));
   OAI22_X1 i_0_0_567 (.A1(n_0_0_471), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_371), 
      .ZN(n_0_0_472));
   OAI22_X1 i_0_0_568 (.A1(n_0_0_472), .A2(i[2]), .B1(n_0_0_23), .B2(n_0_0_428), 
      .ZN(n_0_0_473));
   AOI22_X1 i_0_0_569 (.A1(n_0_0_473), .A2(n_0_0_19), .B1(n_0_0_453), .B2(i[1]), 
      .ZN(n_0_0_474));
   OAI221_X1 i_0_0_570 (.A(n_0_0_100), .B1(i[0]), .B2(n_0_0_474), .C1(n_0_0_15), 
      .C2(n_0_0_464), .ZN(n_0_0_475));
   AOI221_X1 i_0_0_571 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[19]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[3]), .C2(n_0_0_439), .ZN(n_0_0_476));
   OAI22_X1 i_0_0_572 (.A1(n_0_0_476), .A2(i[3]), .B1(n_0_0_9), .B2(n_0_0_378), 
      .ZN(n_0_0_477));
   OAI22_X1 i_0_0_573 (.A1(n_0_0_477), .A2(i[2]), .B1(n_0_0_23), .B2(n_0_0_435), 
      .ZN(n_0_0_478));
   AOI22_X1 i_0_0_574 (.A1(n_0_0_458), .A2(i[1]), .B1(n_0_0_478), .B2(n_0_0_19), 
      .ZN(n_0_0_479));
   OAI22_X1 i_0_0_575 (.A1(n_0_0_479), .A2(i[0]), .B1(n_0_0_469), .B2(n_0_0_15), 
      .ZN(n_0_0_480));
   OAI21_X1 i_0_0_576 (.A(n_0_0_475), .B1(n_0_0_102), .B2(n_0_0_480), .ZN(
      partialProd[35]));
   AOI221_X1 i_0_0_577 (.A(n_0_0_425), .B1(extended_M[4]), .B2(n_0_0_439), 
      .C1(extended_M[20]), .C2(n_0_0_426), .ZN(n_0_0_481));
   OAI22_X1 i_0_0_578 (.A1(n_0_0_481), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_383), 
      .ZN(n_0_0_482));
   AOI22_X1 i_0_0_579 (.A1(n_0_0_23), .A2(n_0_0_482), .B1(n_0_0_442), .B2(i[2]), 
      .ZN(n_0_0_483));
   AOI22_X1 i_0_0_580 (.A1(n_0_0_483), .A2(n_0_0_19), .B1(n_0_0_463), .B2(i[1]), 
      .ZN(n_0_0_484));
   OAI221_X1 i_0_0_581 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_474), .C1(i[0]), 
      .C2(n_0_0_484), .ZN(n_0_0_485));
   AOI221_X1 i_0_0_582 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[4]), .B2(
      n_0_0_439), .C1(extended_M_mul_neg_one[20]), .C2(n_0_0_426), .ZN(n_0_0_486));
   OAI22_X1 i_0_0_583 (.A1(n_0_0_486), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_391), 
      .ZN(n_0_0_487));
   AOI22_X1 i_0_0_584 (.A1(n_0_0_487), .A2(n_0_0_23), .B1(n_0_0_447), .B2(i[2]), 
      .ZN(n_0_0_488));
   OAI22_X1 i_0_0_585 (.A1(n_0_0_488), .A2(i[1]), .B1(n_0_0_468), .B2(n_0_0_19), 
      .ZN(n_0_0_489));
   OAI22_X1 i_0_0_586 (.A1(n_0_0_489), .A2(i[0]), .B1(n_0_0_479), .B2(n_0_0_15), 
      .ZN(n_0_0_490));
   OAI21_X1 i_0_0_587 (.A(n_0_0_485), .B1(n_0_0_102), .B2(n_0_0_490), .ZN(
      partialProd[36]));
   AOI221_X1 i_0_0_588 (.A(n_0_0_425), .B1(extended_M[5]), .B2(n_0_0_439), 
      .C1(extended_M[21]), .C2(n_0_0_426), .ZN(n_0_0_491));
   OAI22_X1 i_0_0_589 (.A1(n_0_0_491), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_397), 
      .ZN(n_0_0_492));
   OAI22_X1 i_0_0_590 (.A1(n_0_0_452), .A2(n_0_0_23), .B1(n_0_0_492), .B2(i[2]), 
      .ZN(n_0_0_493));
   AOI22_X1 i_0_0_591 (.A1(n_0_0_493), .A2(n_0_0_19), .B1(n_0_0_473), .B2(i[1]), 
      .ZN(n_0_0_494));
   OAI221_X1 i_0_0_592 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_484), .C1(i[0]), 
      .C2(n_0_0_494), .ZN(n_0_0_495));
   AOI221_X1 i_0_0_593 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[21]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[5]), .C2(n_0_0_439), .ZN(n_0_0_496));
   OAI22_X1 i_0_0_594 (.A1(n_0_0_496), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_402), 
      .ZN(n_0_0_497));
   OAI22_X1 i_0_0_595 (.A1(n_0_0_497), .A2(i[2]), .B1(n_0_0_457), .B2(n_0_0_23), 
      .ZN(n_0_0_498));
   AOI22_X1 i_0_0_596 (.A1(n_0_0_498), .A2(n_0_0_19), .B1(n_0_0_478), .B2(i[1]), 
      .ZN(n_0_0_499));
   OAI22_X1 i_0_0_597 (.A1(n_0_0_489), .A2(n_0_0_15), .B1(n_0_0_499), .B2(i[0]), 
      .ZN(n_0_0_500));
   OAI21_X1 i_0_0_598 (.A(n_0_0_495), .B1(n_0_0_102), .B2(n_0_0_500), .ZN(
      partialProd[37]));
   AOI221_X1 i_0_0_599 (.A(n_0_0_425), .B1(extended_M[6]), .B2(n_0_0_439), 
      .C1(extended_M[22]), .C2(n_0_0_426), .ZN(n_0_0_501));
   OAI22_X1 i_0_0_600 (.A1(n_0_0_501), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_411), 
      .ZN(n_0_0_502));
   OAI22_X1 i_0_0_601 (.A1(n_0_0_462), .A2(n_0_0_23), .B1(n_0_0_502), .B2(i[2]), 
      .ZN(n_0_0_503));
   AOI22_X1 i_0_0_602 (.A1(n_0_0_19), .A2(n_0_0_503), .B1(n_0_0_483), .B2(i[1]), 
      .ZN(n_0_0_504));
   OAI221_X1 i_0_0_603 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_494), .C1(i[0]), 
      .C2(n_0_0_504), .ZN(n_0_0_505));
   AOI221_X1 i_0_0_604 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[22]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[6]), .C2(n_0_0_439), .ZN(n_0_0_506));
   OAI22_X1 i_0_0_605 (.A1(n_0_0_506), .A2(i[3]), .B1(n_0_0_161), .B2(n_0_0_418), 
      .ZN(n_0_0_507));
   OAI22_X1 i_0_0_606 (.A1(n_0_0_467), .A2(n_0_0_23), .B1(n_0_0_507), .B2(i[2]), 
      .ZN(n_0_0_508));
   OAI22_X1 i_0_0_607 (.A1(n_0_0_508), .A2(i[1]), .B1(n_0_0_488), .B2(n_0_0_19), 
      .ZN(n_0_0_509));
   OAI22_X1 i_0_0_608 (.A1(n_0_0_509), .A2(i[0]), .B1(n_0_0_499), .B2(n_0_0_15), 
      .ZN(n_0_0_510));
   OAI21_X1 i_0_0_609 (.A(n_0_0_505), .B1(n_0_0_102), .B2(n_0_0_510), .ZN(
      partialProd[38]));
   AOI221_X1 i_0_0_610 (.A(n_0_0_425), .B1(extended_M[7]), .B2(n_0_0_439), 
      .C1(extended_M[23]), .C2(n_0_0_426), .ZN(n_0_0_511));
   AOI22_X1 i_0_0_611 (.A1(n_0_0_511), .A2(n_0_0_9), .B1(i[3]), .B2(n_0_0_427), 
      .ZN(n_0_0_512));
   OAI22_X1 i_0_0_612 (.A1(n_0_0_23), .A2(n_0_0_472), .B1(n_0_0_512), .B2(i[2]), 
      .ZN(n_0_0_513));
   AOI22_X1 i_0_0_613 (.A1(i[1]), .A2(n_0_0_493), .B1(n_0_0_513), .B2(n_0_0_19), 
      .ZN(n_0_0_514));
   OAI221_X1 i_0_0_614 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_504), .C1(i[0]), 
      .C2(n_0_0_514), .ZN(n_0_0_515));
   AOI221_X1 i_0_0_615 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[23]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[7]), .C2(n_0_0_439), .ZN(n_0_0_516));
   AOI22_X1 i_0_0_616 (.A1(n_0_0_516), .A2(n_0_0_9), .B1(i[3]), .B2(n_0_0_434), 
      .ZN(n_0_0_517));
   OAI22_X1 i_0_0_617 (.A1(n_0_0_477), .A2(n_0_0_23), .B1(n_0_0_517), .B2(i[2]), 
      .ZN(n_0_0_518));
   AOI22_X1 i_0_0_618 (.A1(i[1]), .A2(n_0_0_498), .B1(n_0_0_518), .B2(n_0_0_19), 
      .ZN(n_0_0_519));
   OAI22_X1 i_0_0_619 (.A1(n_0_0_509), .A2(n_0_0_15), .B1(n_0_0_519), .B2(i[0]), 
      .ZN(n_0_0_520));
   OAI21_X1 i_0_0_620 (.A(n_0_0_515), .B1(n_0_0_102), .B2(n_0_0_520), .ZN(
      partialProd[39]));
   AOI221_X1 i_0_0_621 (.A(n_0_0_425), .B1(extended_M[8]), .B2(n_0_0_439), 
      .C1(extended_M[24]), .C2(n_0_0_426), .ZN(n_0_0_521));
   AOI22_X1 i_0_0_622 (.A1(n_0_0_9), .A2(n_0_0_521), .B1(n_0_0_441), .B2(i[3]), 
      .ZN(n_0_0_522));
   OAI22_X1 i_0_0_623 (.A1(n_0_0_522), .A2(i[2]), .B1(n_0_0_482), .B2(n_0_0_23), 
      .ZN(n_0_0_523));
   AOI22_X1 i_0_0_624 (.A1(n_0_0_523), .A2(n_0_0_19), .B1(n_0_0_503), .B2(i[1]), 
      .ZN(n_0_0_524));
   OAI221_X1 i_0_0_625 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_514), .C1(i[0]), 
      .C2(n_0_0_524), .ZN(n_0_0_525));
   AOI221_X1 i_0_0_626 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[24]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[8]), .C2(n_0_0_439), .ZN(n_0_0_526));
   AOI22_X1 i_0_0_627 (.A1(n_0_0_526), .A2(n_0_0_9), .B1(n_0_0_446), .B2(i[3]), 
      .ZN(n_0_0_527));
   OAI22_X1 i_0_0_628 (.A1(n_0_0_527), .A2(i[2]), .B1(n_0_0_487), .B2(n_0_0_23), 
      .ZN(n_0_0_528));
   AOI22_X1 i_0_0_629 (.A1(n_0_0_528), .A2(n_0_0_19), .B1(n_0_0_508), .B2(i[1]), 
      .ZN(n_0_0_529));
   OAI22_X1 i_0_0_630 (.A1(n_0_0_529), .A2(i[0]), .B1(n_0_0_519), .B2(n_0_0_15), 
      .ZN(n_0_0_530));
   OAI21_X1 i_0_0_631 (.A(n_0_0_525), .B1(n_0_0_102), .B2(n_0_0_530), .ZN(
      partialProd[40]));
   AOI221_X1 i_0_0_632 (.A(n_0_0_425), .B1(extended_M[9]), .B2(n_0_0_439), 
      .C1(extended_M[25]), .C2(n_0_0_426), .ZN(n_0_0_531));
   AOI22_X1 i_0_0_633 (.A1(n_0_0_531), .A2(n_0_0_9), .B1(n_0_0_451), .B2(i[3]), 
      .ZN(n_0_0_532));
   OAI22_X1 i_0_0_634 (.A1(n_0_0_532), .A2(i[2]), .B1(n_0_0_492), .B2(n_0_0_23), 
      .ZN(n_0_0_533));
   AOI22_X1 i_0_0_635 (.A1(n_0_0_533), .A2(n_0_0_19), .B1(n_0_0_513), .B2(i[1]), 
      .ZN(n_0_0_534));
   OAI221_X1 i_0_0_636 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_524), .C1(i[0]), 
      .C2(n_0_0_534), .ZN(n_0_0_535));
   AOI221_X1 i_0_0_637 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[25]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[9]), .C2(n_0_0_439), .ZN(n_0_0_536));
   AOI22_X1 i_0_0_638 (.A1(n_0_0_536), .A2(n_0_0_9), .B1(n_0_0_456), .B2(i[3]), 
      .ZN(n_0_0_537));
   OAI22_X1 i_0_0_639 (.A1(n_0_0_537), .A2(i[2]), .B1(n_0_0_497), .B2(n_0_0_23), 
      .ZN(n_0_0_538));
   AOI22_X1 i_0_0_640 (.A1(n_0_0_538), .A2(n_0_0_19), .B1(n_0_0_518), .B2(i[1]), 
      .ZN(n_0_0_539));
   OAI22_X1 i_0_0_641 (.A1(n_0_0_529), .A2(n_0_0_15), .B1(n_0_0_539), .B2(i[0]), 
      .ZN(n_0_0_540));
   OAI21_X1 i_0_0_642 (.A(n_0_0_535), .B1(n_0_0_102), .B2(n_0_0_540), .ZN(
      partialProd[41]));
   AOI221_X1 i_0_0_643 (.A(n_0_0_425), .B1(extended_M[10]), .B2(n_0_0_439), 
      .C1(extended_M[26]), .C2(n_0_0_426), .ZN(n_0_0_541));
   AOI22_X1 i_0_0_644 (.A1(n_0_0_541), .A2(n_0_0_9), .B1(n_0_0_461), .B2(i[3]), 
      .ZN(n_0_0_542));
   OAI22_X1 i_0_0_645 (.A1(n_0_0_542), .A2(i[2]), .B1(n_0_0_502), .B2(n_0_0_23), 
      .ZN(n_0_0_543));
   AOI22_X1 i_0_0_646 (.A1(n_0_0_19), .A2(n_0_0_543), .B1(n_0_0_523), .B2(i[1]), 
      .ZN(n_0_0_544));
   OAI221_X1 i_0_0_647 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_534), .C1(i[0]), 
      .C2(n_0_0_544), .ZN(n_0_0_545));
   AOI221_X1 i_0_0_648 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[26]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[10]), .C2(n_0_0_439), .ZN(n_0_0_546));
   AOI22_X1 i_0_0_649 (.A1(n_0_0_546), .A2(n_0_0_9), .B1(n_0_0_466), .B2(i[3]), 
      .ZN(n_0_0_547));
   AOI22_X1 i_0_0_650 (.A1(n_0_0_547), .A2(n_0_0_23), .B1(n_0_0_507), .B2(i[2]), 
      .ZN(n_0_0_548));
   AOI22_X1 i_0_0_651 (.A1(n_0_0_548), .A2(n_0_0_19), .B1(n_0_0_528), .B2(i[1]), 
      .ZN(n_0_0_549));
   OAI22_X1 i_0_0_652 (.A1(n_0_0_549), .A2(i[0]), .B1(n_0_0_539), .B2(n_0_0_15), 
      .ZN(n_0_0_550));
   OAI21_X1 i_0_0_653 (.A(n_0_0_545), .B1(n_0_0_102), .B2(n_0_0_550), .ZN(
      partialProd[42]));
   AOI221_X1 i_0_0_654 (.A(n_0_0_425), .B1(extended_M[11]), .B2(n_0_0_439), 
      .C1(extended_M[27]), .C2(n_0_0_426), .ZN(n_0_0_551));
   AOI22_X1 i_0_0_655 (.A1(n_0_0_551), .A2(n_0_0_9), .B1(n_0_0_471), .B2(i[3]), 
      .ZN(n_0_0_552));
   OAI22_X1 i_0_0_656 (.A1(n_0_0_552), .A2(i[2]), .B1(n_0_0_512), .B2(n_0_0_23), 
      .ZN(n_0_0_553));
   AOI22_X1 i_0_0_657 (.A1(i[1]), .A2(n_0_0_533), .B1(n_0_0_553), .B2(n_0_0_19), 
      .ZN(n_0_0_554));
   OAI221_X1 i_0_0_658 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_544), .C1(i[0]), 
      .C2(n_0_0_554), .ZN(n_0_0_555));
   AOI221_X1 i_0_0_659 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[27]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[11]), .C2(n_0_0_439), .ZN(n_0_0_556));
   OAI22_X1 i_0_0_660 (.A1(n_0_0_556), .A2(i[3]), .B1(n_0_0_476), .B2(n_0_0_9), 
      .ZN(n_0_0_557));
   AOI22_X1 i_0_0_661 (.A1(n_0_0_557), .A2(n_0_0_23), .B1(n_0_0_517), .B2(i[2]), 
      .ZN(n_0_0_558));
   OAI22_X1 i_0_0_662 (.A1(n_0_0_538), .A2(n_0_0_19), .B1(n_0_0_558), .B2(i[1]), 
      .ZN(n_0_0_559));
   OAI22_X1 i_0_0_663 (.A1(n_0_0_549), .A2(n_0_0_15), .B1(n_0_0_559), .B2(i[0]), 
      .ZN(n_0_0_560));
   OAI21_X1 i_0_0_664 (.A(n_0_0_555), .B1(n_0_0_102), .B2(n_0_0_560), .ZN(
      partialProd[43]));
   AOI221_X1 i_0_0_665 (.A(n_0_0_425), .B1(extended_M[12]), .B2(n_0_0_439), 
      .C1(extended_M[28]), .C2(n_0_0_426), .ZN(n_0_0_561));
   AOI22_X1 i_0_0_666 (.A1(n_0_0_561), .A2(n_0_0_9), .B1(n_0_0_481), .B2(i[3]), 
      .ZN(n_0_0_562));
   OAI22_X1 i_0_0_667 (.A1(n_0_0_562), .A2(i[2]), .B1(n_0_0_522), .B2(n_0_0_23), 
      .ZN(n_0_0_563));
   AOI22_X1 i_0_0_668 (.A1(n_0_0_563), .A2(n_0_0_19), .B1(n_0_0_543), .B2(i[1]), 
      .ZN(n_0_0_564));
   OAI221_X1 i_0_0_669 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_554), .C1(i[0]), 
      .C2(n_0_0_564), .ZN(n_0_0_565));
   AOI221_X1 i_0_0_670 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[28]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[12]), .C2(n_0_0_439), .ZN(n_0_0_566));
   AOI22_X1 i_0_0_671 (.A1(n_0_0_566), .A2(n_0_0_9), .B1(n_0_0_486), .B2(i[3]), 
      .ZN(n_0_0_567));
   OAI22_X1 i_0_0_672 (.A1(n_0_0_567), .A2(i[2]), .B1(n_0_0_527), .B2(n_0_0_23), 
      .ZN(n_0_0_568));
   AOI22_X1 i_0_0_673 (.A1(n_0_0_548), .A2(i[1]), .B1(n_0_0_568), .B2(n_0_0_19), 
      .ZN(n_0_0_569));
   OAI22_X1 i_0_0_674 (.A1(n_0_0_569), .A2(i[0]), .B1(n_0_0_559), .B2(n_0_0_15), 
      .ZN(n_0_0_570));
   OAI21_X1 i_0_0_675 (.A(n_0_0_565), .B1(n_0_0_102), .B2(n_0_0_570), .ZN(
      partialProd[44]));
   AOI221_X1 i_0_0_676 (.A(n_0_0_425), .B1(extended_M[13]), .B2(n_0_0_439), 
      .C1(extended_M[29]), .C2(n_0_0_426), .ZN(n_0_0_571));
   AOI22_X1 i_0_0_677 (.A1(n_0_0_571), .A2(n_0_0_9), .B1(n_0_0_491), .B2(i[3]), 
      .ZN(n_0_0_572));
   OAI22_X1 i_0_0_678 (.A1(n_0_0_532), .A2(n_0_0_23), .B1(n_0_0_572), .B2(i[2]), 
      .ZN(n_0_0_573));
   AOI22_X1 i_0_0_679 (.A1(n_0_0_573), .A2(n_0_0_19), .B1(n_0_0_553), .B2(i[1]), 
      .ZN(n_0_0_574));
   OAI221_X1 i_0_0_680 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_564), .C1(i[0]), 
      .C2(n_0_0_574), .ZN(n_0_0_575));
   AOI221_X1 i_0_0_681 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[29]), .B2(
      n_0_0_426), .C1(extended_M_mul_neg_one[13]), .C2(n_0_0_439), .ZN(n_0_0_576));
   AOI22_X1 i_0_0_682 (.A1(n_0_0_576), .A2(n_0_0_9), .B1(n_0_0_496), .B2(i[3]), 
      .ZN(n_0_0_577));
   OAI22_X1 i_0_0_683 (.A1(n_0_0_537), .A2(n_0_0_23), .B1(n_0_0_577), .B2(i[2]), 
      .ZN(n_0_0_578));
   OAI22_X1 i_0_0_684 (.A1(n_0_0_578), .A2(i[1]), .B1(n_0_0_558), .B2(n_0_0_19), 
      .ZN(n_0_0_579));
   OAI22_X1 i_0_0_685 (.A1(n_0_0_579), .A2(i[0]), .B1(n_0_0_569), .B2(n_0_0_15), 
      .ZN(n_0_0_580));
   OAI21_X1 i_0_0_686 (.A(n_0_0_575), .B1(n_0_0_102), .B2(n_0_0_580), .ZN(
      partialProd[45]));
   AOI221_X1 i_0_0_687 (.A(n_0_0_425), .B1(extended_M[14]), .B2(n_0_0_439), 
      .C1(extended_M[30]), .C2(n_0_0_426), .ZN(n_0_0_581));
   AOI22_X1 i_0_0_688 (.A1(n_0_0_581), .A2(n_0_0_9), .B1(n_0_0_501), .B2(i[3]), 
      .ZN(n_0_0_582));
   OAI22_X1 i_0_0_689 (.A1(n_0_0_542), .A2(n_0_0_23), .B1(n_0_0_582), .B2(i[2]), 
      .ZN(n_0_0_583));
   AOI22_X1 i_0_0_690 (.A1(n_0_0_19), .A2(n_0_0_583), .B1(n_0_0_563), .B2(i[1]), 
      .ZN(n_0_0_584));
   OAI221_X1 i_0_0_691 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_574), .C1(i[0]), 
      .C2(n_0_0_584), .ZN(n_0_0_585));
   AOI221_X1 i_0_0_692 (.A(n_0_0_433), .B1(extended_M_mul_neg_one[14]), .B2(
      n_0_0_439), .C1(extended_M_mul_neg_one[30]), .C2(n_0_0_426), .ZN(n_0_0_586));
   AOI22_X1 i_0_0_693 (.A1(n_0_0_586), .A2(n_0_0_9), .B1(n_0_0_506), .B2(i[3]), 
      .ZN(n_0_0_587));
   OAI22_X1 i_0_0_694 (.A1(n_0_0_587), .A2(i[2]), .B1(n_0_0_547), .B2(n_0_0_23), 
      .ZN(n_0_0_588));
   AOI22_X1 i_0_0_695 (.A1(n_0_0_588), .A2(n_0_0_19), .B1(n_0_0_568), .B2(i[1]), 
      .ZN(n_0_0_589));
   OAI22_X1 i_0_0_696 (.A1(n_0_0_579), .A2(n_0_0_15), .B1(n_0_0_589), .B2(i[0]), 
      .ZN(n_0_0_590));
   OAI21_X1 i_0_0_697 (.A(n_0_0_585), .B1(n_0_0_102), .B2(n_0_0_590), .ZN(
      partialProd[46]));
   INV_X1 i_0_0_698 (.A(n_0_0_424), .ZN(n_0_0_591));
   AOI21_X1 i_0_0_699 (.A(n_0_0_591), .B1(n_0_0_439), .B2(extended_M[15]), 
      .ZN(n_0_0_592));
   AOI22_X1 i_0_0_700 (.A1(n_0_0_511), .A2(i[3]), .B1(n_0_0_9), .B2(n_0_0_592), 
      .ZN(n_0_0_593));
   OAI22_X1 i_0_0_701 (.A1(n_0_0_552), .A2(n_0_0_23), .B1(n_0_0_593), .B2(i[2]), 
      .ZN(n_0_0_594));
   AOI22_X1 i_0_0_702 (.A1(n_0_0_573), .A2(i[1]), .B1(n_0_0_594), .B2(n_0_0_19), 
      .ZN(n_0_0_595));
   OAI221_X1 i_0_0_703 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_584), .C1(i[0]), 
      .C2(n_0_0_595), .ZN(n_0_0_596));
   INV_X1 i_0_0_704 (.A(n_0_0_432), .ZN(n_0_0_597));
   AOI21_X1 i_0_0_705 (.A(n_0_0_597), .B1(n_0_0_439), .B2(
      extended_M_mul_neg_one[15]), .ZN(n_0_0_598));
   AOI22_X1 i_0_0_706 (.A1(n_0_0_516), .A2(i[3]), .B1(n_0_0_9), .B2(n_0_0_598), 
      .ZN(n_0_0_599));
   OAI22_X1 i_0_0_707 (.A1(n_0_0_557), .A2(n_0_0_23), .B1(n_0_0_599), .B2(i[2]), 
      .ZN(n_0_0_600));
   AOI22_X1 i_0_0_708 (.A1(n_0_0_578), .A2(i[1]), .B1(n_0_0_600), .B2(n_0_0_19), 
      .ZN(n_0_0_601));
   OAI22_X1 i_0_0_709 (.A1(n_0_0_589), .A2(n_0_0_15), .B1(n_0_0_601), .B2(i[0]), 
      .ZN(n_0_0_602));
   OAI21_X1 i_0_0_710 (.A(n_0_0_596), .B1(n_0_0_102), .B2(n_0_0_602), .ZN(
      partialProd[47]));
   NOR2_X1 i_0_0_711 (.A1(n_0_0_591), .A2(i[3]), .ZN(n_0_0_603));
   INV_X1 i_0_0_712 (.A(n_0_0_603), .ZN(n_0_0_604));
   AOI21_X1 i_0_0_713 (.A(n_0_0_604), .B1(n_0_0_253), .B2(i[5]), .ZN(n_0_0_605));
   AOI21_X1 i_0_0_714 (.A(n_0_0_605), .B1(n_0_0_521), .B2(i[3]), .ZN(n_0_0_606));
   OAI22_X1 i_0_0_715 (.A1(n_0_0_562), .A2(n_0_0_23), .B1(n_0_0_606), .B2(i[2]), 
      .ZN(n_0_0_607));
   AOI22_X1 i_0_0_716 (.A1(n_0_0_583), .A2(i[1]), .B1(n_0_0_607), .B2(n_0_0_19), 
      .ZN(n_0_0_608));
   OAI221_X1 i_0_0_717 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_595), .C1(i[0]), 
      .C2(n_0_0_608), .ZN(n_0_0_609));
   AOI21_X1 i_0_0_718 (.A(n_0_0_597), .B1(n_0_0_260), .B2(i[5]), .ZN(n_0_0_610));
   AOI22_X1 i_0_0_719 (.A1(n_0_0_526), .A2(i[3]), .B1(n_0_0_610), .B2(n_0_0_9), 
      .ZN(n_0_0_611));
   AOI22_X1 i_0_0_720 (.A1(n_0_0_567), .A2(i[2]), .B1(n_0_0_611), .B2(n_0_0_23), 
      .ZN(n_0_0_612));
   AOI22_X1 i_0_0_721 (.A1(n_0_0_588), .A2(i[1]), .B1(n_0_0_612), .B2(n_0_0_19), 
      .ZN(n_0_0_613));
   OAI22_X1 i_0_0_722 (.A1(n_0_0_613), .A2(i[0]), .B1(n_0_0_601), .B2(n_0_0_15), 
      .ZN(n_0_0_614));
   OAI21_X1 i_0_0_723 (.A(n_0_0_609), .B1(n_0_0_102), .B2(n_0_0_614), .ZN(
      partialProd[48]));
   INV_X1 i_0_0_724 (.A(n_0_0_266), .ZN(n_0_0_615));
   AOI21_X1 i_0_0_725 (.A(n_0_0_604), .B1(n_0_0_615), .B2(i[5]), .ZN(n_0_0_616));
   AOI21_X1 i_0_0_726 (.A(n_0_0_616), .B1(n_0_0_531), .B2(i[3]), .ZN(n_0_0_617));
   OAI22_X1 i_0_0_727 (.A1(n_0_0_572), .A2(n_0_0_23), .B1(n_0_0_617), .B2(i[2]), 
      .ZN(n_0_0_618));
   AOI22_X1 i_0_0_728 (.A1(n_0_0_594), .A2(i[1]), .B1(n_0_0_618), .B2(n_0_0_19), 
      .ZN(n_0_0_619));
   OAI221_X1 i_0_0_729 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_608), .C1(i[0]), 
      .C2(n_0_0_619), .ZN(n_0_0_620));
   AOI21_X1 i_0_0_730 (.A(n_0_0_597), .B1(n_0_0_272), .B2(i[5]), .ZN(n_0_0_621));
   AOI22_X1 i_0_0_731 (.A1(n_0_0_536), .A2(i[3]), .B1(n_0_0_9), .B2(n_0_0_621), 
      .ZN(n_0_0_622));
   OAI22_X1 i_0_0_732 (.A1(n_0_0_577), .A2(n_0_0_23), .B1(n_0_0_622), .B2(i[2]), 
      .ZN(n_0_0_623));
   AOI22_X1 i_0_0_733 (.A1(n_0_0_623), .A2(n_0_0_19), .B1(n_0_0_600), .B2(i[1]), 
      .ZN(n_0_0_624));
   OAI22_X1 i_0_0_734 (.A1(n_0_0_613), .A2(n_0_0_15), .B1(n_0_0_624), .B2(i[0]), 
      .ZN(n_0_0_625));
   OAI21_X1 i_0_0_735 (.A(n_0_0_620), .B1(n_0_0_102), .B2(n_0_0_625), .ZN(
      partialProd[49]));
   INV_X1 i_0_0_736 (.A(n_0_0_278), .ZN(n_0_0_626));
   AOI21_X1 i_0_0_737 (.A(n_0_0_591), .B1(n_0_0_626), .B2(i[5]), .ZN(n_0_0_627));
   AOI22_X1 i_0_0_738 (.A1(n_0_0_541), .A2(i[3]), .B1(n_0_0_627), .B2(n_0_0_9), 
      .ZN(n_0_0_628));
   OAI22_X1 i_0_0_739 (.A1(n_0_0_582), .A2(n_0_0_23), .B1(n_0_0_628), .B2(i[2]), 
      .ZN(n_0_0_629));
   AOI22_X1 i_0_0_740 (.A1(n_0_0_629), .A2(n_0_0_19), .B1(n_0_0_607), .B2(i[1]), 
      .ZN(n_0_0_630));
   OAI221_X1 i_0_0_741 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_619), .C1(i[0]), 
      .C2(n_0_0_630), .ZN(n_0_0_631));
   INV_X1 i_0_0_742 (.A(n_0_0_283), .ZN(n_0_0_632));
   AOI21_X1 i_0_0_743 (.A(n_0_0_597), .B1(n_0_0_632), .B2(i[5]), .ZN(n_0_0_633));
   AOI22_X1 i_0_0_744 (.A1(n_0_0_546), .A2(i[3]), .B1(n_0_0_9), .B2(n_0_0_633), 
      .ZN(n_0_0_634));
   OAI22_X1 i_0_0_745 (.A1(n_0_0_587), .A2(n_0_0_23), .B1(n_0_0_634), .B2(i[2]), 
      .ZN(n_0_0_635));
   AOI22_X1 i_0_0_746 (.A1(n_0_0_612), .A2(i[1]), .B1(n_0_0_635), .B2(n_0_0_19), 
      .ZN(n_0_0_636));
   OAI22_X1 i_0_0_747 (.A1(n_0_0_636), .A2(i[0]), .B1(n_0_0_624), .B2(n_0_0_15), 
      .ZN(n_0_0_637));
   OAI21_X1 i_0_0_748 (.A(n_0_0_631), .B1(n_0_0_102), .B2(n_0_0_637), .ZN(
      partialProd[50]));
   INV_X1 i_0_0_749 (.A(n_0_0_288), .ZN(n_0_0_638));
   AOI21_X1 i_0_0_750 (.A(n_0_0_604), .B1(n_0_0_638), .B2(i[5]), .ZN(n_0_0_639));
   AOI21_X1 i_0_0_751 (.A(n_0_0_639), .B1(n_0_0_551), .B2(i[3]), .ZN(n_0_0_640));
   OAI22_X1 i_0_0_752 (.A1(n_0_0_593), .A2(n_0_0_23), .B1(n_0_0_640), .B2(i[2]), 
      .ZN(n_0_0_641));
   AOI22_X1 i_0_0_753 (.A1(n_0_0_618), .A2(i[1]), .B1(n_0_0_641), .B2(n_0_0_19), 
      .ZN(n_0_0_642));
   OAI221_X1 i_0_0_754 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_630), .C1(i[0]), 
      .C2(n_0_0_642), .ZN(n_0_0_643));
   INV_X1 i_0_0_755 (.A(n_0_0_293), .ZN(n_0_0_644));
   AOI21_X1 i_0_0_756 (.A(n_0_0_597), .B1(n_0_0_644), .B2(i[5]), .ZN(n_0_0_645));
   AOI22_X1 i_0_0_757 (.A1(n_0_0_556), .A2(i[3]), .B1(n_0_0_9), .B2(n_0_0_645), 
      .ZN(n_0_0_646));
   OAI22_X1 i_0_0_758 (.A1(n_0_0_599), .A2(n_0_0_23), .B1(n_0_0_646), .B2(i[2]), 
      .ZN(n_0_0_647));
   AOI22_X1 i_0_0_759 (.A1(n_0_0_623), .A2(i[1]), .B1(n_0_0_647), .B2(n_0_0_19), 
      .ZN(n_0_0_648));
   OAI22_X1 i_0_0_760 (.A1(n_0_0_636), .A2(n_0_0_15), .B1(n_0_0_648), .B2(i[0]), 
      .ZN(n_0_0_649));
   OAI21_X1 i_0_0_761 (.A(n_0_0_643), .B1(n_0_0_102), .B2(n_0_0_649), .ZN(
      partialProd[51]));
   AOI21_X1 i_0_0_762 (.A(n_0_0_604), .B1(n_0_0_385), .B2(i[5]), .ZN(n_0_0_650));
   AOI21_X1 i_0_0_763 (.A(n_0_0_650), .B1(n_0_0_561), .B2(i[3]), .ZN(n_0_0_651));
   OAI22_X1 i_0_0_764 (.A1(n_0_0_651), .A2(i[2]), .B1(n_0_0_606), .B2(n_0_0_23), 
      .ZN(n_0_0_652));
   AOI22_X1 i_0_0_765 (.A1(n_0_0_629), .A2(i[1]), .B1(n_0_0_652), .B2(n_0_0_19), 
      .ZN(n_0_0_653));
   OAI221_X1 i_0_0_766 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_642), .C1(i[0]), 
      .C2(n_0_0_653), .ZN(n_0_0_654));
   NAND2_X1 i_0_0_767 (.A1(n_0_0_432), .A2(n_0_0_9), .ZN(n_0_0_655));
   INV_X1 i_0_0_768 (.A(n_0_0_303), .ZN(n_0_0_656));
   AOI21_X1 i_0_0_769 (.A(n_0_0_655), .B1(n_0_0_656), .B2(i[5]), .ZN(n_0_0_657));
   AOI21_X1 i_0_0_770 (.A(n_0_0_657), .B1(n_0_0_566), .B2(i[3]), .ZN(n_0_0_658));
   OAI22_X1 i_0_0_771 (.A1(n_0_0_611), .A2(n_0_0_23), .B1(n_0_0_658), .B2(i[2]), 
      .ZN(n_0_0_659));
   AOI22_X1 i_0_0_772 (.A1(n_0_0_635), .A2(i[1]), .B1(n_0_0_659), .B2(n_0_0_19), 
      .ZN(n_0_0_660));
   OAI22_X1 i_0_0_773 (.A1(n_0_0_648), .A2(n_0_0_15), .B1(n_0_0_660), .B2(i[0]), 
      .ZN(n_0_0_661));
   OAI21_X1 i_0_0_774 (.A(n_0_0_654), .B1(n_0_0_102), .B2(n_0_0_661), .ZN(
      partialProd[52]));
   INV_X1 i_0_0_775 (.A(n_0_0_308), .ZN(n_0_0_662));
   AOI21_X1 i_0_0_776 (.A(n_0_0_604), .B1(n_0_0_662), .B2(i[5]), .ZN(n_0_0_663));
   AOI21_X1 i_0_0_777 (.A(n_0_0_663), .B1(n_0_0_571), .B2(i[3]), .ZN(n_0_0_664));
   OAI22_X1 i_0_0_778 (.A1(n_0_0_617), .A2(n_0_0_23), .B1(n_0_0_664), .B2(i[2]), 
      .ZN(n_0_0_665));
   AOI22_X1 i_0_0_779 (.A1(n_0_0_641), .A2(i[1]), .B1(n_0_0_665), .B2(n_0_0_19), 
      .ZN(n_0_0_666));
   OAI221_X1 i_0_0_780 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_653), .C1(i[0]), 
      .C2(n_0_0_666), .ZN(n_0_0_667));
   AOI21_X1 i_0_0_781 (.A(n_0_0_655), .B1(n_0_0_404), .B2(i[5]), .ZN(n_0_0_668));
   AOI21_X1 i_0_0_782 (.A(n_0_0_668), .B1(n_0_0_576), .B2(i[3]), .ZN(n_0_0_669));
   OAI22_X1 i_0_0_783 (.A1(n_0_0_622), .A2(n_0_0_23), .B1(n_0_0_669), .B2(i[2]), 
      .ZN(n_0_0_670));
   AOI22_X1 i_0_0_784 (.A1(i[1]), .A2(n_0_0_647), .B1(n_0_0_670), .B2(n_0_0_19), 
      .ZN(n_0_0_671));
   OAI22_X1 i_0_0_785 (.A1(n_0_0_660), .A2(n_0_0_15), .B1(n_0_0_671), .B2(i[0]), 
      .ZN(n_0_0_672));
   OAI21_X1 i_0_0_786 (.A(n_0_0_667), .B1(n_0_0_102), .B2(n_0_0_672), .ZN(
      partialProd[53]));
   AOI21_X1 i_0_0_787 (.A(n_0_0_604), .B1(n_0_0_410), .B2(i[5]), .ZN(n_0_0_673));
   AOI21_X1 i_0_0_788 (.A(n_0_0_673), .B1(n_0_0_581), .B2(i[3]), .ZN(n_0_0_674));
   OAI22_X1 i_0_0_789 (.A1(n_0_0_628), .A2(n_0_0_23), .B1(n_0_0_674), .B2(i[2]), 
      .ZN(n_0_0_675));
   AOI22_X1 i_0_0_790 (.A1(n_0_0_675), .A2(n_0_0_19), .B1(n_0_0_652), .B2(i[1]), 
      .ZN(n_0_0_676));
   OAI221_X1 i_0_0_791 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_666), .C1(i[0]), 
      .C2(n_0_0_676), .ZN(n_0_0_677));
   INV_X1 i_0_0_792 (.A(n_0_0_323), .ZN(n_0_0_678));
   AOI21_X1 i_0_0_793 (.A(n_0_0_655), .B1(n_0_0_678), .B2(i[5]), .ZN(n_0_0_679));
   AOI21_X1 i_0_0_794 (.A(n_0_0_679), .B1(n_0_0_586), .B2(i[3]), .ZN(n_0_0_680));
   OAI22_X1 i_0_0_795 (.A1(n_0_0_634), .A2(n_0_0_23), .B1(n_0_0_680), .B2(i[2]), 
      .ZN(n_0_0_681));
   AOI22_X1 i_0_0_796 (.A1(n_0_0_659), .A2(i[1]), .B1(n_0_0_681), .B2(n_0_0_19), 
      .ZN(n_0_0_682));
   OAI22_X1 i_0_0_797 (.A1(n_0_0_682), .A2(i[0]), .B1(n_0_0_671), .B2(n_0_0_15), 
      .ZN(n_0_0_683));
   OAI21_X1 i_0_0_798 (.A(n_0_0_677), .B1(n_0_0_102), .B2(n_0_0_683), .ZN(
      partialProd[54]));
   OR2_X1 i_0_0_799 (.A1(n_0_0_328), .A2(n_0_0_10), .ZN(n_0_0_684));
   AOI22_X1 i_0_0_800 (.A1(n_0_0_684), .A2(n_0_0_603), .B1(n_0_0_592), .B2(i[3]), 
      .ZN(n_0_0_685));
   OAI22_X1 i_0_0_801 (.A1(n_0_0_640), .A2(n_0_0_23), .B1(i[2]), .B2(n_0_0_685), 
      .ZN(n_0_0_686));
   AOI22_X1 i_0_0_802 (.A1(n_0_0_665), .A2(i[1]), .B1(n_0_0_686), .B2(n_0_0_19), 
      .ZN(n_0_0_687));
   OAI221_X1 i_0_0_803 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_676), .C1(i[0]), 
      .C2(n_0_0_687), .ZN(n_0_0_688));
   INV_X1 i_0_0_804 (.A(extended_M_mul_neg_one[63]), .ZN(n_0_0_689));
   OAI21_X1 i_0_0_805 (.A(n_0_0_97), .B1(n_0_0_689), .B2(i[3]), .ZN(n_0_0_690));
   INV_X1 i_0_0_806 (.A(n_0_0_333), .ZN(n_0_0_691));
   OAI21_X1 i_0_0_807 (.A(n_0_0_690), .B1(n_0_0_691), .B2(n_0_0_10), .ZN(
      n_0_0_692));
   OAI21_X1 i_0_0_808 (.A(n_0_0_692), .B1(n_0_0_9), .B2(n_0_0_598), .ZN(
      n_0_0_693));
   OAI22_X1 i_0_0_809 (.A1(n_0_0_646), .A2(n_0_0_23), .B1(i[2]), .B2(n_0_0_693), 
      .ZN(n_0_0_694));
   AOI22_X1 i_0_0_810 (.A1(n_0_0_670), .A2(i[1]), .B1(n_0_0_694), .B2(n_0_0_19), 
      .ZN(n_0_0_695));
   OAI22_X1 i_0_0_811 (.A1(n_0_0_682), .A2(n_0_0_15), .B1(n_0_0_695), .B2(i[0]), 
      .ZN(n_0_0_696));
   OAI21_X1 i_0_0_812 (.A(n_0_0_688), .B1(n_0_0_102), .B2(n_0_0_696), .ZN(
      partialProd[55]));
   INV_X1 i_0_0_813 (.A(n_0_0_340), .ZN(n_0_0_697));
   AOI21_X1 i_0_0_814 (.A(n_0_0_591), .B1(n_0_0_697), .B2(i[5]), .ZN(n_0_0_698));
   INV_X1 i_0_0_815 (.A(n_0_0_698), .ZN(n_0_0_699));
   OAI22_X1 i_0_0_816 (.A1(n_0_0_651), .A2(n_0_0_23), .B1(n_0_0_699), .B2(i[2]), 
      .ZN(n_0_0_700));
   AOI22_X1 i_0_0_817 (.A1(n_0_0_675), .A2(i[1]), .B1(n_0_0_700), .B2(n_0_0_19), 
      .ZN(n_0_0_701));
   OAI221_X1 i_0_0_818 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_687), .C1(i[0]), 
      .C2(n_0_0_701), .ZN(n_0_0_702));
   INV_X1 i_0_0_819 (.A(n_0_0_610), .ZN(n_0_0_703));
   NAND2_X1 i_0_0_820 (.A1(n_0_0_345), .A2(i[5]), .ZN(n_0_0_704));
   AOI22_X1 i_0_0_821 (.A1(n_0_0_703), .A2(i[3]), .B1(n_0_0_704), .B2(n_0_0_690), 
      .ZN(n_0_0_705));
   INV_X1 i_0_0_822 (.A(n_0_0_705), .ZN(n_0_0_706));
   OAI22_X1 i_0_0_823 (.A1(n_0_0_658), .A2(n_0_0_23), .B1(n_0_0_706), .B2(i[2]), 
      .ZN(n_0_0_707));
   AOI22_X1 i_0_0_824 (.A1(n_0_0_681), .A2(i[1]), .B1(n_0_0_707), .B2(n_0_0_19), 
      .ZN(n_0_0_708));
   OAI22_X1 i_0_0_825 (.A1(n_0_0_695), .A2(n_0_0_15), .B1(n_0_0_708), .B2(i[0]), 
      .ZN(n_0_0_709));
   OAI21_X1 i_0_0_826 (.A(n_0_0_702), .B1(n_0_0_102), .B2(n_0_0_709), .ZN(
      partialProd[56]));
   NOR2_X1 i_0_0_827 (.A1(extended_M[63]), .A2(i[5]), .ZN(n_0_0_710));
   NOR3_X1 i_0_0_828 (.A1(n_0_0_615), .A2(n_0_0_9), .A3(n_0_0_10), .ZN(n_0_0_711));
   INV_X1 i_0_0_829 (.A(n_0_0_97), .ZN(n_0_0_712));
   AOI211_X1 i_0_0_830 (.A(n_0_0_710), .B(n_0_0_711), .C1(n_0_0_712), .C2(
      n_0_0_350), .ZN(n_0_0_713));
   OAI22_X1 i_0_0_831 (.A1(n_0_0_664), .A2(n_0_0_23), .B1(n_0_0_713), .B2(i[2]), 
      .ZN(n_0_0_714));
   AOI22_X1 i_0_0_832 (.A1(n_0_0_714), .A2(n_0_0_19), .B1(n_0_0_686), .B2(i[1]), 
      .ZN(n_0_0_715));
   OAI221_X1 i_0_0_833 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_701), .C1(i[0]), 
      .C2(n_0_0_715), .ZN(n_0_0_716));
   INV_X1 i_0_0_834 (.A(n_0_0_355), .ZN(n_0_0_717));
   OAI21_X1 i_0_0_835 (.A(n_0_0_690), .B1(n_0_0_717), .B2(n_0_0_10), .ZN(
      n_0_0_718));
   OAI21_X1 i_0_0_836 (.A(n_0_0_718), .B1(n_0_0_621), .B2(n_0_0_9), .ZN(
      n_0_0_719));
   OAI22_X1 i_0_0_837 (.A1(n_0_0_669), .A2(n_0_0_23), .B1(n_0_0_719), .B2(i[2]), 
      .ZN(n_0_0_720));
   AOI22_X1 i_0_0_838 (.A1(i[1]), .A2(n_0_0_694), .B1(n_0_0_720), .B2(n_0_0_19), 
      .ZN(n_0_0_721));
   OAI22_X1 i_0_0_839 (.A1(n_0_0_708), .A2(n_0_0_15), .B1(n_0_0_721), .B2(i[0]), 
      .ZN(n_0_0_722));
   OAI21_X1 i_0_0_840 (.A(n_0_0_716), .B1(n_0_0_102), .B2(n_0_0_722), .ZN(
      partialProd[57]));
   OR2_X1 i_0_0_841 (.A1(n_0_0_360), .A2(n_0_0_10), .ZN(n_0_0_723));
   AOI22_X1 i_0_0_842 (.A1(n_0_0_627), .A2(i[3]), .B1(n_0_0_723), .B2(n_0_0_603), 
      .ZN(n_0_0_724));
   OAI22_X1 i_0_0_843 (.A1(n_0_0_674), .A2(n_0_0_23), .B1(i[2]), .B2(n_0_0_724), 
      .ZN(n_0_0_725));
   AOI22_X1 i_0_0_844 (.A1(n_0_0_700), .A2(i[1]), .B1(n_0_0_725), .B2(n_0_0_19), 
      .ZN(n_0_0_726));
   OAI221_X1 i_0_0_845 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_715), .C1(i[0]), 
      .C2(n_0_0_726), .ZN(n_0_0_727));
   INV_X1 i_0_0_846 (.A(n_0_0_633), .ZN(n_0_0_728));
   NAND2_X1 i_0_0_847 (.A1(n_0_0_365), .A2(i[5]), .ZN(n_0_0_729));
   AOI22_X1 i_0_0_848 (.A1(n_0_0_728), .A2(i[3]), .B1(n_0_0_729), .B2(n_0_0_690), 
      .ZN(n_0_0_730));
   INV_X1 i_0_0_849 (.A(n_0_0_730), .ZN(n_0_0_731));
   OAI22_X1 i_0_0_850 (.A1(n_0_0_680), .A2(n_0_0_23), .B1(n_0_0_731), .B2(i[2]), 
      .ZN(n_0_0_732));
   AOI22_X1 i_0_0_851 (.A1(n_0_0_732), .A2(n_0_0_19), .B1(n_0_0_707), .B2(i[1]), 
      .ZN(n_0_0_733));
   OAI22_X1 i_0_0_852 (.A1(n_0_0_721), .A2(n_0_0_15), .B1(n_0_0_733), .B2(i[0]), 
      .ZN(n_0_0_734));
   OAI21_X1 i_0_0_853 (.A(n_0_0_727), .B1(n_0_0_102), .B2(n_0_0_734), .ZN(
      partialProd[58]));
   NAND3_X1 i_0_0_854 (.A1(n_0_0_288), .A2(i[3]), .A3(i[5]), .ZN(n_0_0_735));
   INV_X1 i_0_0_855 (.A(n_0_0_710), .ZN(n_0_0_736));
   INV_X1 i_0_0_856 (.A(n_0_0_371), .ZN(n_0_0_737));
   OAI211_X1 i_0_0_857 (.A(n_0_0_735), .B(n_0_0_736), .C1(n_0_0_97), .C2(
      n_0_0_737), .ZN(n_0_0_738));
   INV_X1 i_0_0_858 (.A(n_0_0_738), .ZN(n_0_0_739));
   AOI22_X1 i_0_0_859 (.A1(n_0_0_739), .A2(n_0_0_23), .B1(i[2]), .B2(n_0_0_685), 
      .ZN(n_0_0_740));
   AOI22_X1 i_0_0_860 (.A1(n_0_0_714), .A2(i[1]), .B1(n_0_0_740), .B2(n_0_0_19), 
      .ZN(n_0_0_741));
   OAI221_X1 i_0_0_861 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_726), .C1(i[0]), 
      .C2(n_0_0_741), .ZN(n_0_0_742));
   OAI21_X1 i_0_0_862 (.A(n_0_0_690), .B1(n_0_0_377), .B2(n_0_0_10), .ZN(
      n_0_0_743));
   OAI21_X1 i_0_0_863 (.A(n_0_0_743), .B1(n_0_0_645), .B2(n_0_0_9), .ZN(
      n_0_0_744));
   OAI22_X1 i_0_0_864 (.A1(n_0_0_744), .A2(i[2]), .B1(n_0_0_693), .B2(n_0_0_23), 
      .ZN(n_0_0_745));
   AOI22_X1 i_0_0_865 (.A1(n_0_0_720), .A2(i[1]), .B1(n_0_0_19), .B2(n_0_0_745), 
      .ZN(n_0_0_746));
   OAI22_X1 i_0_0_866 (.A1(n_0_0_733), .A2(n_0_0_15), .B1(n_0_0_746), .B2(i[0]), 
      .ZN(n_0_0_747));
   OAI21_X1 i_0_0_867 (.A(n_0_0_742), .B1(n_0_0_102), .B2(n_0_0_747), .ZN(
      partialProd[59]));
   INV_X1 i_0_0_868 (.A(n_0_0_386), .ZN(n_0_0_748));
   AOI21_X1 i_0_0_869 (.A(n_0_0_591), .B1(n_0_0_748), .B2(i[5]), .ZN(n_0_0_749));
   AOI222_X1 i_0_0_870 (.A1(n_0_0_725), .A2(i[1]), .B1(n_0_0_698), .B2(n_0_0_21), 
      .C1(n_0_0_749), .C2(n_0_0_13), .ZN(n_0_0_750));
   OAI221_X1 i_0_0_871 (.A(n_0_0_100), .B1(n_0_0_15), .B2(n_0_0_741), .C1(i[0]), 
      .C2(n_0_0_750), .ZN(n_0_0_751));
   AOI21_X1 i_0_0_872 (.A(n_0_0_597), .B1(n_0_0_392), .B2(i[5]), .ZN(n_0_0_752));
   AOI222_X1 i_0_0_873 (.A1(n_0_0_732), .A2(i[1]), .B1(n_0_0_705), .B2(n_0_0_21), 
      .C1(n_0_0_13), .C2(n_0_0_752), .ZN(n_0_0_753));
   OAI22_X1 i_0_0_874 (.A1(n_0_0_753), .A2(i[0]), .B1(n_0_0_746), .B2(n_0_0_15), 
      .ZN(n_0_0_754));
   OAI21_X1 i_0_0_875 (.A(n_0_0_751), .B1(n_0_0_102), .B2(n_0_0_754), .ZN(
      partialProd[60]));
   NOR3_X1 i_0_0_876 (.A1(n_0_0_662), .A2(n_0_0_9), .A3(n_0_0_10), .ZN(n_0_0_755));
   AOI211_X1 i_0_0_877 (.A(n_0_0_710), .B(n_0_0_755), .C1(n_0_0_712), .C2(
      n_0_0_397), .ZN(n_0_0_756));
   AOI22_X1 i_0_0_878 (.A1(n_0_0_756), .A2(n_0_0_23), .B1(n_0_0_713), .B2(i[2]), 
      .ZN(n_0_0_757));
   AOI22_X1 i_0_0_879 (.A1(n_0_0_757), .A2(n_0_0_19), .B1(n_0_0_740), .B2(i[1]), 
      .ZN(n_0_0_758));
   OAI221_X1 i_0_0_880 (.A(n_0_0_100), .B1(i[0]), .B2(n_0_0_758), .C1(n_0_0_15), 
      .C2(n_0_0_750), .ZN(n_0_0_759));
   OAI211_X1 i_0_0_881 (.A(n_0_0_13), .B(n_0_0_432), .C1(n_0_0_405), .C2(
      n_0_0_10), .ZN(n_0_0_760));
   OAI21_X1 i_0_0_882 (.A(n_0_0_760), .B1(n_0_0_20), .B2(n_0_0_719), .ZN(
      n_0_0_761));
   AOI21_X1 i_0_0_883 (.A(n_0_0_761), .B1(n_0_0_745), .B2(i[1]), .ZN(n_0_0_762));
   OAI22_X1 i_0_0_884 (.A1(n_0_0_753), .A2(n_0_0_15), .B1(i[0]), .B2(n_0_0_762), 
      .ZN(n_0_0_763));
   OAI21_X1 i_0_0_885 (.A(n_0_0_759), .B1(n_0_0_102), .B2(n_0_0_763), .ZN(
      partialProd[61]));
   AOI22_X1 i_0_0_886 (.A1(n_0_0_705), .A2(n_0_0_18), .B1(n_0_0_21), .B2(
      n_0_0_730), .ZN(n_0_0_764));
   AOI21_X1 i_0_0_887 (.A(n_0_0_597), .B1(n_0_0_419), .B2(i[5]), .ZN(n_0_0_765));
   AOI22_X1 i_0_0_888 (.A1(n_0_0_765), .A2(n_0_0_13), .B1(n_0_0_752), .B2(
      n_0_0_25), .ZN(n_0_0_766));
   NAND3_X1 i_0_0_889 (.A1(n_0_0_764), .A2(n_0_0_766), .A3(n_0_0_15), .ZN(
      n_0_0_767));
   INV_X1 i_0_0_890 (.A(n_0_0_762), .ZN(n_0_0_768));
   OAI21_X1 i_0_0_891 (.A(n_0_0_767), .B1(n_0_0_768), .B2(n_0_0_15), .ZN(
      n_0_0_769));
   NAND2_X1 i_0_0_892 (.A1(n_0_0_107), .A2(n_0_0_769), .ZN(n_0_0_770));
   AOI21_X1 i_0_0_893 (.A(n_0_0_710), .B1(n_0_0_413), .B2(i[5]), .ZN(n_0_0_771));
   OAI22_X1 i_0_0_894 (.A1(n_0_0_771), .A2(n_0_0_34), .B1(n_0_0_724), .B2(
      n_0_0_20), .ZN(n_0_0_772));
   AOI221_X1 i_0_0_895 (.A(n_0_0_772), .B1(n_0_0_25), .B2(n_0_0_749), .C1(
      n_0_0_18), .C2(n_0_0_698), .ZN(n_0_0_773));
   AOI22_X1 i_0_0_896 (.A1(n_0_0_758), .A2(i[0]), .B1(n_0_0_773), .B2(n_0_0_15), 
      .ZN(n_0_0_774));
   OAI21_X1 i_0_0_897 (.A(n_0_0_770), .B1(n_0_0_101), .B2(n_0_0_774), .ZN(
      partialProd[62]));
   AOI221_X1 i_0_0_898 (.A(i[0]), .B1(n_0_0_21), .B2(n_0_0_738), .C1(n_0_0_757), 
      .C2(i[1]), .ZN(n_0_0_775));
   NAND2_X1 i_0_0_899 (.A1(i[4]), .A2(i[5]), .ZN(n_0_0_776));
   INV_X1 i_0_0_900 (.A(n_0_0_776), .ZN(n_0_0_777));
   OAI221_X1 i_0_0_901 (.A(n_0_0_9), .B1(n_0_0_776), .B2(extended_M[15]), 
      .C1(n_0_0_777), .C2(extended_M[63]), .ZN(n_0_0_778));
   INV_X1 i_0_0_902 (.A(n_0_0_684), .ZN(n_0_0_779));
   OAI21_X1 i_0_0_903 (.A(i[3]), .B1(n_0_0_779), .B2(n_0_0_591), .ZN(n_0_0_780));
   NAND3_X1 i_0_0_904 (.A1(n_0_0_778), .A2(n_0_0_780), .A3(n_0_0_13), .ZN(
      n_0_0_781));
   AOI22_X1 i_0_0_905 (.A1(n_0_0_775), .A2(n_0_0_781), .B1(n_0_0_773), .B2(i[0]), 
      .ZN(n_0_0_782));
   OAI21_X1 i_0_0_906 (.A(n_0_0_770), .B1(n_0_0_101), .B2(n_0_0_782), .ZN(
      partialProd[63]));
   AND2_X1 i_0_0_907 (.A1(n_0_0_8), .A2(n_0_0_4), .ZN(n_0_163));
   AND2_X1 i_0_0_908 (.A1(n_0_0_8), .A2(n_0_0_5), .ZN(n_0_164));
   AND2_X1 i_0_0_909 (.A1(n_0_0_8), .A2(n_0_0_6), .ZN(n_0_165));
   AND2_X1 i_0_0_910 (.A1(n_0_0_8), .A2(n_0_0_7), .ZN(n_0_166));
   INV_X1 i_0_0_911 (.A(n_0_0_3), .ZN(n_0_0_783));
   AOI221_X1 i_0_0_912 (.A(start), .B1(i[5]), .B2(n_0_0_3), .C1(n_0_0_10), 
      .C2(n_0_0_783), .ZN(n_0_167));
   NOR2_X1 i_0_0_913 (.A1(i[0]), .A2(start), .ZN(n_0_162));
   AND2_X1 i_0_0_914 (.A1(n_0_0_98), .A2(n_0_162), .ZN(n_0_169));
   INV_X1 i_0_0_915 (.A(n_0_169), .ZN(n_0_168));
   DFF_X1 \Acc_reg[63]  (.D(n_0_161), .CK(n_0_1), .Q(Acc[63]), .QN());
   DFF_X1 \Acc_reg[62]  (.D(n_0_160), .CK(n_0_1), .Q(Acc[62]), .QN());
   DFF_X1 \Acc_reg[61]  (.D(n_0_159), .CK(n_0_1), .Q(Acc[61]), .QN());
   DFF_X1 \Acc_reg[60]  (.D(n_0_158), .CK(n_0_1), .Q(Acc[60]), .QN());
   DFF_X1 \Acc_reg[59]  (.D(n_0_157), .CK(n_0_1), .Q(Acc[59]), .QN());
   DFF_X1 \Acc_reg[58]  (.D(n_0_156), .CK(n_0_1), .Q(Acc[58]), .QN());
   DFF_X1 \Acc_reg[57]  (.D(n_0_155), .CK(n_0_1), .Q(Acc[57]), .QN());
   DFF_X1 \Acc_reg[56]  (.D(n_0_154), .CK(n_0_1), .Q(Acc[56]), .QN());
   DFF_X1 \Acc_reg[55]  (.D(n_0_153), .CK(n_0_1), .Q(Acc[55]), .QN());
   DFF_X1 \Acc_reg[54]  (.D(n_0_152), .CK(n_0_1), .Q(Acc[54]), .QN());
   DFF_X1 \Acc_reg[53]  (.D(n_0_151), .CK(n_0_1), .Q(Acc[53]), .QN());
   DFF_X1 \Acc_reg[52]  (.D(n_0_150), .CK(n_0_1), .Q(Acc[52]), .QN());
   DFF_X1 \Acc_reg[51]  (.D(n_0_149), .CK(n_0_1), .Q(Acc[51]), .QN());
   DFF_X1 \Acc_reg[50]  (.D(n_0_148), .CK(n_0_1), .Q(Acc[50]), .QN());
   DFF_X1 \Acc_reg[49]  (.D(n_0_147), .CK(n_0_1), .Q(Acc[49]), .QN());
   DFF_X1 \Acc_reg[48]  (.D(n_0_146), .CK(n_0_1), .Q(Acc[48]), .QN());
   DFF_X1 \Acc_reg[47]  (.D(n_0_145), .CK(n_0_1), .Q(Acc[47]), .QN());
   DFF_X1 \Acc_reg[46]  (.D(n_0_144), .CK(n_0_1), .Q(Acc[46]), .QN());
   DFF_X1 \Acc_reg[45]  (.D(n_0_143), .CK(n_0_1), .Q(Acc[45]), .QN());
   DFF_X1 \Acc_reg[44]  (.D(n_0_142), .CK(n_0_1), .Q(Acc[44]), .QN());
   DFF_X1 \Acc_reg[43]  (.D(n_0_141), .CK(n_0_1), .Q(Acc[43]), .QN());
   DFF_X1 \Acc_reg[42]  (.D(n_0_140), .CK(n_0_1), .Q(Acc[42]), .QN());
   DFF_X1 \Acc_reg[41]  (.D(n_0_139), .CK(n_0_1), .Q(Acc[41]), .QN());
   DFF_X1 \Acc_reg[40]  (.D(n_0_138), .CK(n_0_1), .Q(Acc[40]), .QN());
   DFF_X1 \Acc_reg[39]  (.D(n_0_137), .CK(n_0_1), .Q(Acc[39]), .QN());
   DFF_X1 \Acc_reg[38]  (.D(n_0_136), .CK(n_0_1), .Q(Acc[38]), .QN());
   DFF_X1 \Acc_reg[37]  (.D(n_0_135), .CK(n_0_1), .Q(Acc[37]), .QN());
   DFF_X1 \Acc_reg[36]  (.D(n_0_134), .CK(n_0_1), .Q(Acc[36]), .QN());
   DFF_X1 \Acc_reg[35]  (.D(n_0_133), .CK(n_0_1), .Q(Acc[35]), .QN());
   DFF_X1 \Acc_reg[34]  (.D(n_0_132), .CK(n_0_1), .Q(Acc[34]), .QN());
   DFF_X1 \Acc_reg[33]  (.D(n_0_131), .CK(n_0_1), .Q(Acc[33]), .QN());
   DFF_X1 \Acc_reg[32]  (.D(n_0_130), .CK(n_0_1), .Q(Acc[32]), .QN());
   DFF_X1 \Acc_reg[31]  (.D(n_0_129), .CK(n_0_1), .Q(Acc[31]), .QN());
   DFF_X1 \Acc_reg[30]  (.D(n_0_128), .CK(n_0_1), .Q(Acc[30]), .QN());
   DFF_X1 \Acc_reg[29]  (.D(n_0_127), .CK(n_0_1), .Q(Acc[29]), .QN());
   DFF_X1 \Acc_reg[28]  (.D(n_0_126), .CK(n_0_1), .Q(Acc[28]), .QN());
   DFF_X1 \Acc_reg[27]  (.D(n_0_125), .CK(n_0_1), .Q(Acc[27]), .QN());
   DFF_X1 \Acc_reg[26]  (.D(n_0_124), .CK(n_0_1), .Q(Acc[26]), .QN());
   DFF_X1 \Acc_reg[25]  (.D(n_0_123), .CK(n_0_1), .Q(Acc[25]), .QN());
   DFF_X1 \Acc_reg[24]  (.D(n_0_122), .CK(n_0_1), .Q(Acc[24]), .QN());
   DFF_X1 \Acc_reg[23]  (.D(n_0_121), .CK(n_0_1), .Q(Acc[23]), .QN());
   DFF_X1 \Acc_reg[22]  (.D(n_0_120), .CK(n_0_1), .Q(Acc[22]), .QN());
   DFF_X1 \Acc_reg[21]  (.D(n_0_119), .CK(n_0_1), .Q(Acc[21]), .QN());
   DFF_X1 \Acc_reg[20]  (.D(n_0_118), .CK(n_0_1), .Q(Acc[20]), .QN());
   DFF_X1 \Acc_reg[19]  (.D(n_0_117), .CK(n_0_1), .Q(Acc[19]), .QN());
   DFF_X1 \Acc_reg[18]  (.D(n_0_116), .CK(n_0_1), .Q(Acc[18]), .QN());
   DFF_X1 \Acc_reg[17]  (.D(n_0_115), .CK(n_0_1), .Q(Acc[17]), .QN());
   DFF_X1 \Acc_reg[16]  (.D(n_0_114), .CK(n_0_1), .Q(Acc[16]), .QN());
   DFF_X1 \Acc_reg[15]  (.D(n_0_113), .CK(n_0_1), .Q(Acc[15]), .QN());
   DFF_X1 \Acc_reg[14]  (.D(n_0_112), .CK(n_0_1), .Q(Acc[14]), .QN());
   DFF_X1 \Acc_reg[13]  (.D(n_0_111), .CK(n_0_1), .Q(Acc[13]), .QN());
   DFF_X1 \Acc_reg[12]  (.D(n_0_110), .CK(n_0_1), .Q(Acc[12]), .QN());
   DFF_X1 \Acc_reg[11]  (.D(n_0_109), .CK(n_0_1), .Q(Acc[11]), .QN());
   DFF_X1 \Acc_reg[10]  (.D(n_0_108), .CK(n_0_1), .Q(Acc[10]), .QN());
   DFF_X1 \Acc_reg[9]  (.D(n_0_107), .CK(n_0_1), .Q(Acc[9]), .QN());
   DFF_X1 \Acc_reg[8]  (.D(n_0_106), .CK(n_0_1), .Q(Acc[8]), .QN());
   DFF_X1 \Acc_reg[7]  (.D(n_0_105), .CK(n_0_1), .Q(Acc[7]), .QN());
   DFF_X1 \Acc_reg[6]  (.D(n_0_104), .CK(n_0_1), .Q(Acc[6]), .QN());
   DFF_X1 \Acc_reg[5]  (.D(n_0_103), .CK(n_0_1), .Q(Acc[5]), .QN());
   DFF_X1 \Acc_reg[4]  (.D(n_0_102), .CK(n_0_1), .Q(Acc[4]), .QN());
   DFF_X1 \Acc_reg[3]  (.D(n_0_101), .CK(n_0_1), .Q(Acc[3]), .QN());
   DFF_X1 \Acc_reg[2]  (.D(n_0_100), .CK(n_0_1), .Q(Acc[2]), .QN());
   DFF_X1 \Acc_reg[1]  (.D(n_0_99), .CK(n_0_1), .Q(Acc[1]), .QN());
   DFF_X1 \Acc_reg[0]  (.D(n_0_98), .CK(n_0_1), .Q(Acc[0]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[63]  (.D(n_0_32), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[63]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[30]  (.D(n_0_31), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[30]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[29]  (.D(n_0_30), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[29]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[28]  (.D(n_0_29), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[28]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[27]  (.D(n_0_28), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[27]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[26]  (.D(n_0_27), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[26]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[25]  (.D(n_0_26), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[25]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[24]  (.D(n_0_25), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[24]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[23]  (.D(n_0_24), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[23]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[22]  (.D(n_0_23), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[22]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[21]  (.D(n_0_22), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[21]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[20]  (.D(n_0_21), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[20]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[19]  (.D(n_0_20), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[19]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[18]  (.D(n_0_19), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[18]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[17]  (.D(n_0_18), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[17]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[16]  (.D(n_0_17), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[16]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[15]  (.D(n_0_16), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[15]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[14]  (.D(n_0_15), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[14]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[13]  (.D(n_0_14), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[13]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[12]  (.D(n_0_13), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[12]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[11]  (.D(n_0_12), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[11]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[10]  (.D(n_0_11), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[10]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[9]  (.D(n_0_10), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[9]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[8]  (.D(n_0_9), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[8]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[7]  (.D(n_0_8), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[7]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[6]  (.D(n_0_7), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[6]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[5]  (.D(n_0_6), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[5]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[4]  (.D(n_0_5), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[4]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[3]  (.D(n_0_4), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[3]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[2]  (.D(n_0_3), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[2]), .QN());
   DFF_X1 \extended_M_mul_neg_one_reg[1]  (.D(n_0_2), .CK(n_0_33), .Q(
      extended_M_mul_neg_one[1]), .QN());
   DFF_X1 \i_reg[5]  (.D(n_0_167), .CK(n_0_1), .Q(i[5]), .QN());
   DFF_X1 \i_reg[4]  (.D(n_0_166), .CK(n_0_1), .Q(i[4]), .QN());
   DFF_X1 \i_reg[3]  (.D(n_0_165), .CK(n_0_1), .Q(i[3]), .QN());
   DFF_X1 \i_reg[2]  (.D(n_0_164), .CK(n_0_1), .Q(i[2]), .QN());
   DFF_X1 \i_reg[1]  (.D(n_0_163), .CK(n_0_1), .Q(i[1]), .QN());
   DFF_X1 \i_reg[0]  (.D(n_0_162), .CK(n_0_1), .Q(i[0]), .QN());
   DFF_X1 \extended_M_reg[63]  (.D(A_reg[31]), .CK(n_0_33), .Q(extended_M[63]), 
      .QN());
   DFF_X1 \extended_M_reg[30]  (.D(A_reg[30]), .CK(n_0_33), .Q(extended_M[30]), 
      .QN());
   DFF_X1 \extended_M_reg[29]  (.D(A_reg[29]), .CK(n_0_33), .Q(extended_M[29]), 
      .QN());
   DFF_X1 \extended_M_reg[28]  (.D(A_reg[28]), .CK(n_0_33), .Q(extended_M[28]), 
      .QN());
   DFF_X1 \extended_M_reg[27]  (.D(A_reg[27]), .CK(n_0_33), .Q(extended_M[27]), 
      .QN());
   DFF_X1 \extended_M_reg[26]  (.D(A_reg[26]), .CK(n_0_33), .Q(extended_M[26]), 
      .QN());
   DFF_X1 \extended_M_reg[25]  (.D(A_reg[25]), .CK(n_0_33), .Q(extended_M[25]), 
      .QN());
   DFF_X1 \extended_M_reg[24]  (.D(A_reg[24]), .CK(n_0_33), .Q(extended_M[24]), 
      .QN());
   DFF_X1 \extended_M_reg[23]  (.D(A_reg[23]), .CK(n_0_33), .Q(extended_M[23]), 
      .QN());
   DFF_X1 \extended_M_reg[22]  (.D(A_reg[22]), .CK(n_0_33), .Q(extended_M[22]), 
      .QN());
   DFF_X1 \extended_M_reg[21]  (.D(A_reg[21]), .CK(n_0_33), .Q(extended_M[21]), 
      .QN());
   DFF_X1 \extended_M_reg[20]  (.D(A_reg[20]), .CK(n_0_33), .Q(extended_M[20]), 
      .QN());
   DFF_X1 \extended_M_reg[19]  (.D(A_reg[19]), .CK(n_0_33), .Q(extended_M[19]), 
      .QN());
   DFF_X1 \extended_M_reg[18]  (.D(A_reg[18]), .CK(n_0_33), .Q(extended_M[18]), 
      .QN());
   DFF_X1 \extended_M_reg[17]  (.D(A_reg[17]), .CK(n_0_33), .Q(extended_M[17]), 
      .QN());
   DFF_X1 \extended_M_reg[16]  (.D(A_reg[16]), .CK(n_0_33), .Q(extended_M[16]), 
      .QN());
   DFF_X1 \extended_M_reg[15]  (.D(A_reg[15]), .CK(n_0_33), .Q(extended_M[15]), 
      .QN());
   DFF_X1 \extended_M_reg[14]  (.D(A_reg[14]), .CK(n_0_33), .Q(extended_M[14]), 
      .QN());
   DFF_X1 \extended_M_reg[13]  (.D(A_reg[13]), .CK(n_0_33), .Q(extended_M[13]), 
      .QN());
   DFF_X1 \extended_M_reg[12]  (.D(A_reg[12]), .CK(n_0_33), .Q(extended_M[12]), 
      .QN());
   DFF_X1 \extended_M_reg[11]  (.D(A_reg[11]), .CK(n_0_33), .Q(extended_M[11]), 
      .QN());
   DFF_X1 \extended_M_reg[10]  (.D(A_reg[10]), .CK(n_0_33), .Q(extended_M[10]), 
      .QN());
   DFF_X1 \extended_M_reg[9]  (.D(A_reg[9]), .CK(n_0_33), .Q(extended_M[9]), 
      .QN());
   DFF_X1 \extended_M_reg[8]  (.D(A_reg[8]), .CK(n_0_33), .Q(extended_M[8]), 
      .QN());
   DFF_X1 \extended_M_reg[7]  (.D(A_reg[7]), .CK(n_0_33), .Q(extended_M[7]), 
      .QN());
   DFF_X1 \extended_M_reg[6]  (.D(A_reg[6]), .CK(n_0_33), .Q(extended_M[6]), 
      .QN());
   DFF_X1 \extended_M_reg[5]  (.D(A_reg[5]), .CK(n_0_33), .Q(extended_M[5]), 
      .QN());
   DFF_X1 \extended_M_reg[4]  (.D(A_reg[4]), .CK(n_0_33), .Q(extended_M[4]), 
      .QN());
   DFF_X1 \extended_M_reg[3]  (.D(A_reg[3]), .CK(n_0_33), .Q(extended_M[3]), 
      .QN());
   DFF_X1 \extended_M_reg[2]  (.D(A_reg[2]), .CK(n_0_33), .Q(extended_M[2]), 
      .QN());
   DFF_X1 \extended_M_reg[1]  (.D(A_reg[1]), .CK(n_0_33), .Q(extended_M[1]), 
      .QN());
   DFF_X1 \Q_reg[32]  (.D(B_reg[31]), .CK(n_0_33), .Q(Q[32]), .QN());
   DFF_X1 \Q_reg[31]  (.D(B_reg[30]), .CK(n_0_33), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(B_reg[29]), .CK(n_0_33), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(B_reg[28]), .CK(n_0_33), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(B_reg[27]), .CK(n_0_33), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(B_reg[26]), .CK(n_0_33), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(B_reg[25]), .CK(n_0_33), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(B_reg[24]), .CK(n_0_33), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(B_reg[23]), .CK(n_0_33), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(B_reg[22]), .CK(n_0_33), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(B_reg[21]), .CK(n_0_33), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(B_reg[20]), .CK(n_0_33), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(B_reg[19]), .CK(n_0_33), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(B_reg[18]), .CK(n_0_33), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(B_reg[17]), .CK(n_0_33), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(B_reg[16]), .CK(n_0_33), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(B_reg[15]), .CK(n_0_33), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(B_reg[14]), .CK(n_0_33), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(B_reg[13]), .CK(n_0_33), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(B_reg[12]), .CK(n_0_33), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(B_reg[11]), .CK(n_0_33), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(B_reg[10]), .CK(n_0_33), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(B_reg[9]), .CK(n_0_33), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(B_reg[8]), .CK(n_0_33), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(B_reg[7]), .CK(n_0_33), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(B_reg[6]), .CK(n_0_33), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(B_reg[5]), .CK(n_0_33), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(B_reg[4]), .CK(n_0_33), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(B_reg[3]), .CK(n_0_33), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(B_reg[2]), .CK(n_0_33), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(B_reg[1]), .CK(n_0_33), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(B_reg[0]), .CK(n_0_33), .Q(Q[1]), .QN());
   CLKGATETST_X1 clk_gate_Acc_reg (.CK(clk), .E(n_0_168), .SE(1'b0), .GCK(n_0_1));
   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(start), .SE(1'b0), .GCK(n_0_33));
   DFF_X1 \extended_M_reg[0]  (.D(A_reg[0]), .CK(n_0_33), .Q(extended_M[0]), 
      .QN());
endmodule
